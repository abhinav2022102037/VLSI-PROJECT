magic
tech scmos
timestamp 1699599481
<< metal1 >>
rect 15 95 33 98
rect 15 47 18 95
rect 26 72 34 76
rect 55 73 58 76
rect 26 58 30 72
rect 58 58 66 61
rect 26 54 30 56
rect -4 21 -2 25
rect 63 4 66 58
rect 75 20 77 25
rect 48 1 66 4
<< m2contact >>
rect 55 20 60 25
rect 69 20 75 25
<< metal2 >>
rect 60 21 69 24
use not  not_0
timestamp 1698566035
transform 1 0 33 0 1 79
box 0 -21 25 19
use NAND  NAND_0
timestamp 1699598546
transform 1 0 -1 0 1 28
box -1 -27 57 30
<< labels >>
rlabel metal1 55 73 58 76 1 out
rlabel metal1 -4 21 -2 25 3 in1
rlabel metal1 75 20 77 25 7 in2
rlabel metal1 48 1 66 4 1 gnd
rlabel metal1 15 95 20 98 5 vdd
<< end >>
