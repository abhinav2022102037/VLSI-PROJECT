ALU circuit
.include TSMC_180nm.txt
.include AND.sub
.include NAND.sub
.include NOT.sub
.include XOR.sub
.include comparator.sub
.include OR.sub
.include NOR.sub
.include XNOR.sub
.include 3inputAND.sub
.include 4inputAND.sub
.include 5inputAND.sub
.include 4inputOR.sub
.include 3inputOR.sub
.include addersubtractor.sub
.include andblock.sub
.include enable.sub
.include fulladder.sub
.include twotofourdecoder.sub
.include ALU.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}
.global gnd

Vdd node_x gnd 'SUPPLY'
V_in_A3 node_A3 gnd PULSE(1.8 0 0ns 100ps 100ps 20ns 70ns)
V_in_A2 node_A2 gnd PULSE(0 1.8 0ns 100ps 100ps 70ns 100ns)
V_in_A1 node_A1 gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 80ns)
V_in_A0 node_A0 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_B3 node_B3 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 80ns)
V_in_B2 node_B2 gnd PULSE(1.8 0 0ns 100ps 100ps 70ns 110ns)
V_in_B1 node_B1 gnd PULSE(0 1.8 0ns 100ps 100ps 30ns 90ns)
V_in_B0 node_B0 gnd PULSE(1.8 0 0ns 100ps 100ps 50ns 70ns)
V_in_S1 S1 gnd 0
V_in_S0 S0 gnd 1.8



X1000 S0 S1 node_A3 node_A2 node_A1 node_A0 node_B3 node_B2 node_B1 node_B0 adder3 adder2 adder1 adder0 carry equal lesser greater and3 and2 and1 and0 node_x gnd ALU
C3 adder3 gnd 3.5f
C2 adder2 gnd 3.5f
C1 adder1 gnd 3.5f
C0 adder0 gnd 3.5f
C4 carry gnd 3.5f
C5 and3 gnd 3.5f
C6 and2 gnd 3.5f
C7 and1 gnd 3.5f
C8 and0 gnd 3.5f
C9 equal gnd 3.5f
C10 greater gnd 3.5f
C11 lesser gnd 3.5f
.tran 1n 400n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(node_A0) v(node_A1)+2 v(node_A2)+4 v(node_A3)+6 v(node_B0)+8 v(node_B1)+10 v(node_B2)+12 v(node_B3)+14
plot v(S0) v(S1)+2 v(adder0)+4 v(adder1)+6 v(adder2)+8 v(adder3)+10 v(carry)+12
plot v(S0) v(S1)+2 v(lesser)+4 v(equal)+6 v(greater)+8 
plot v(S0) v(S1)+2 v(and0)+4 v(and1)+6 v(and2)+8 v(and3)+10 
.end
.endc


