XNOR gate
.include TSMC_180nm.txt
.include NOT.sub
.include XOR.sub
.include XNOR.sub
.include NAND.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}
.global gnd

Vdd node_x gnd 'SUPPLY'
V_in_a node_a gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b node_b gnd PULSE(0 1.8 0ns 100ps 100ps 30ns 70ns)

X17 node_a node_b node_out node_x gnd XNOR
.tran 1n 200n

.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(node_a) v(node_b)+2 v(node_out)+4
hardcopy XNOR.ps v(node_a) v(node_b)+2 v(node_out)+4
.end
.endc


