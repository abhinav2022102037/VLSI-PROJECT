magic
tech scmos
timestamp 1699603457
<< metal1 >>
rect -119 132 -116 165
rect -36 133 -33 161
rect 54 135 57 165
rect 151 138 154 166
rect 142 135 154 138
rect -133 129 -115 132
rect -44 130 -33 133
rect 46 132 57 135
rect -25 81 -16 84
rect 65 83 81 86
rect 162 83 165 86
rect -114 78 -106 81
rect -195 0 -192 77
rect -128 6 -125 52
rect -105 21 -102 78
rect -25 54 -22 81
rect 65 58 68 83
rect 62 55 68 58
rect -25 51 45 54
rect 30 40 46 43
rect 71 40 144 43
rect -105 18 6 21
rect 161 21 164 83
rect 168 45 171 160
rect 45 17 47 21
rect 63 18 164 21
rect -128 3 6 6
rect 30 3 47 6
rect 80 0 83 18
rect -195 -3 83 0
rect -19 -5 -15 -3
rect -133 -14 -128 -12
rect -105 -13 -100 -11
<< m2contact >>
rect -133 151 -128 156
rect -92 152 -87 157
rect -44 152 -39 157
rect -2 152 3 157
rect 46 154 51 159
rect 95 155 100 160
rect 143 157 148 162
rect 163 156 168 161
rect -129 52 -124 57
rect -133 5 -128 10
rect -96 52 -90 58
rect -36 56 -31 62
rect 54 63 59 68
rect -11 58 -6 63
rect 57 54 62 59
rect 86 60 91 66
rect 40 46 45 51
rect 144 39 149 44
rect -105 13 -100 18
rect 27 17 32 22
rect 40 17 45 22
rect 167 40 172 45
rect -133 -12 -128 -7
rect -105 -11 -100 -6
<< metal2 >>
rect -128 153 -92 156
rect -39 153 -2 156
rect 51 155 95 158
rect 148 158 163 161
rect 59 66 91 67
rect 59 64 86 66
rect -124 52 -96 55
rect -31 59 -11 62
rect 32 55 57 58
rect 32 18 35 55
rect 41 22 44 46
rect 149 40 167 43
rect -132 -7 -129 5
rect -104 -6 -101 13
use AND  AND_3
timestamp 1699599481
transform 1 0 -191 0 1 56
box -4 1 77 98
use AND  AND_2
timestamp 1699599481
transform 1 0 85 0 1 62
box -4 1 77 98
use AND  AND_1
timestamp 1699599481
transform 1 0 -12 0 1 59
box -4 1 77 98
use AND  AND_0
timestamp 1699599481
transform 1 0 -102 0 1 57
box -4 1 77 98
use not  not_1
timestamp 1698566035
transform 1 0 46 0 1 24
box 0 -21 25 19
use not  not_0
timestamp 1698566035
transform 1 0 5 0 1 24
box 0 -21 25 19
<< labels >>
rlabel metal1 -36 159 -33 161 5 D1
rlabel metal1 54 161 57 165 5 D0
rlabel metal1 -119 160 -116 165 5 D3
rlabel metal1 -133 -14 -128 -12 1 gnd
rlabel metal1 -105 -13 -100 -11 1 S0
rlabel metal1 -19 -5 -15 -3 1 S1
rlabel metal1 151 163 154 166 5 D2
rlabel metal1 168 155 171 160 7 vdd
<< end >>
