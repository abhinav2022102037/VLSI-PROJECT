enable circuit
.include TSMC_180nm.txt
.include AND.sub
.include NAND.sub
.include NOT.sub
.include enable.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}
.global gnd

Vdd node_x gnd 'SUPPLY'
V_in_A3 node_A3 gnd PULSE(0 1.8 0ns 100ps 100ps 80ns 160ns)
V_in_A2 node_A2 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_A1 node_A1 gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 80ns)
V_in_A0 node_A0 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_B3 node_B3 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_B2 node_B2 gnd PULSE(0 1.8 0ns 100ps 100ps 80ns 160ns)
V_in_B1 node_B1 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_B0 node_B0 gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 80ns)
V_in_enable En gnd  PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
X24 En node_A3 node_A2 node_A1 node_A0 node_B3 node_B2 node_B1 node_B0 A_out3 A_out2 A_out1 A_out0 B_out3 B_out2 B_out1 B_out0 node_x gnd enable

.tran 1n 300n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(En)-2 v(node_A0) v(node_A1)+2 v(node_A2)+4 v(node_A3)+6 v(node_B0)+8 v(node_B1)+10 v(node_B2)+12 v(node_B3)+14 v(A_out0)+16 v(A_out1)+18 v(A_out2)+20 v(A_out3)+22 v(B_out0)+24 v(B_out1)+26 v(B_out2)+28 v(B_out3)+30 
.end
.endc


