ALU
.include TSMC_180nm.txt
.option scale=0.09u
.param SUPPLY = 1.8
.param LAMBDA = 0.09u

.param width_P = 8*LAMBDA
.param width_N = 4*LAMBDA

.global vdd

Vdd vdd gnd 'SUPPLY'
V_in_A3 A3 gnd PULSE(1.8 0 0ns 100ps 100ps 30ns 70ns)
V_in_A2 A2 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 100ns)
V_in_A1 A1 gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 80ns)
V_in_A0 A0 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_B3 B3 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 90ns)
V_in_B2 B2 gnd PULSE(1.8 0 0ns 100ps 100ps 70ns 110ns)
V_in_B1 B1 gnd PULSE(0 1.8 0ns 100ps 100ps 30ns 90ns)
V_in_B0 B0 gnd PULSE(1.8 0 0ns 100ps 100ps 50ns 80ns)
V_in_S1 S1 gnd 0
V_in_S0 S0 gnd 1.8

M1000 addersubtractor_0/fulladder_0/AND_0/not_0/in addersubtractor_0/XOR_0/out addersubtractor_0/fulladder_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1001 addersubtractor_0/fulladder_0/AND_0/not_0/in addersubtractor_0/XOR_0/out vdd vdd CMOSP w=4 l=2
+  ad=40 pd=36 as=6270 ps=5638
M1002 gnd enableblock_0/A_out3 addersubtractor_0/fulladder_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=3920 pd=3528 as=0 ps=0
M1003 vdd enableblock_0/A_out3 addersubtractor_0/fulladder_0/AND_0/not_0/in addersubtractor_0/fulladder_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1005 addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/AND_0/not_0/in vdd addersubtractor_0/fulladder_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1006 addersubtractor_0/fulladder_0/AND_1/not_0/in S0 addersubtractor_0/fulladder_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1007 addersubtractor_0/fulladder_0/AND_1/not_0/in S0 vdd addersubtractor_0/fulladder_0/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1008 gnd addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 vdd addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/AND_1/not_0/in addersubtractor_0/fulladder_0/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 addersubtractor_0/fulladder_0/OR_0/in1 addersubtractor_0/fulladder_0/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1011 addersubtractor_0/fulladder_0/OR_0/in1 addersubtractor_0/fulladder_0/AND_1/not_0/in vdd addersubtractor_0/fulladder_0/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1012 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 enableblock_0/A_out3 addersubtractor_0/fulladder_0/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1013 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 enableblock_0/A_out3 vdd addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1014 gnd addersubtractor_0/XOR_0/out addersubtractor_0/fulladder_0/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 vdd addersubtractor_0/XOR_0/out addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 enableblock_0/A_out3 addersubtractor_0/fulladder_0/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1017 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 enableblock_0/A_out3 vdd addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1018 gnd addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 vdd addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1021 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 vdd addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1022 gnd addersubtractor_0/XOR_0/out addersubtractor_0/fulladder_0/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 vdd addersubtractor_0/XOR_0/out addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1025 addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 vdd addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1026 gnd addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 vdd addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_0/OR_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1029 addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_0/OR_0/NOT_0/in vdd addersubtractor_0/fulladder_0/OR_0/NOT_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1030 addersubtractor_0/fulladder_0/OR_0/NOT_0/in addersubtractor_0/fulladder_0/OR_0/in1 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1031 addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_0/OR_0/in1 vdd addersubtractor_0/fulladder_0/OR_0/NOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1032 gnd addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/OR_0/NOT_0/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1033 addersubtractor_0/fulladder_0/OR_0/NOT_0/in addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_0/OR_0/NOR_0/w_32_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1034 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 S0 addersubtractor_0/fulladder_0/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1035 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 S0 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1036 gnd addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 vdd addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 S0 addersubtractor_0/fulladder_0/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1039 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 S0 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1040 gnd addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1043 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1044 gnd addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1045 vdd addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 adder0 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1047 adder0 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1048 gnd addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1049 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 adder0 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/XOR_1/out addersubtractor_0/fulladder_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1051 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/XOR_1/out vdd addersubtractor_0/fulladder_1/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1052 gnd enableblock_0/A_out1 addersubtractor_0/fulladder_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1053 vdd enableblock_0/A_out1 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/fulladder_1/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 addersubtractor_0/fulladder_1/OR_0/in2 addersubtractor_0/fulladder_1/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1055 addersubtractor_0/fulladder_1/OR_0/in2 addersubtractor_0/fulladder_1/AND_0/not_0/in vdd addersubtractor_0/fulladder_1/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1056 addersubtractor_0/fulladder_1/AND_1/not_0/in addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1057 addersubtractor_0/fulladder_1/AND_1/not_0/in addersubtractor_0/fulladder_0/C vdd addersubtractor_0/fulladder_1/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1058 gnd addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1059 vdd addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/AND_1/not_0/in addersubtractor_0/fulladder_1/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 addersubtractor_0/fulladder_1/OR_0/in1 addersubtractor_0/fulladder_1/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1061 addersubtractor_0/fulladder_1/OR_0/in1 addersubtractor_0/fulladder_1/AND_1/not_0/in vdd addersubtractor_0/fulladder_1/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1062 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 enableblock_0/A_out1 addersubtractor_0/fulladder_1/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1063 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 enableblock_0/A_out1 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1064 gnd addersubtractor_0/XOR_1/out addersubtractor_0/fulladder_1/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 vdd addersubtractor_0/XOR_1/out addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 enableblock_0/A_out1 addersubtractor_0/fulladder_1/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1067 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 enableblock_0/A_out1 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1068 gnd addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1069 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1071 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1072 gnd addersubtractor_0/XOR_1/out addersubtractor_0/fulladder_1/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 vdd addersubtractor_0/XOR_1/out addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1075 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1076 gnd addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_1/OR_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1079 addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_1/OR_0/NOT_0/in vdd addersubtractor_0/fulladder_1/OR_0/NOT_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1080 addersubtractor_0/fulladder_1/OR_0/NOT_0/in addersubtractor_0/fulladder_1/OR_0/in1 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1081 addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_1/OR_0/in1 vdd addersubtractor_0/fulladder_1/OR_0/NOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1082 gnd addersubtractor_0/fulladder_1/OR_0/in2 addersubtractor_0/fulladder_1/OR_0/NOT_0/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 addersubtractor_0/fulladder_1/OR_0/NOT_0/in addersubtractor_0/fulladder_1/OR_0/in2 addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_1/OR_0/NOR_0/w_32_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1084 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_1/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1085 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/C vdd addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1086 gnd addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 vdd addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_1/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1089 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_0/C vdd addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1090 gnd addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1092 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1093 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1094 gnd addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 vdd addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 adder1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1097 adder1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1098 gnd addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 adder1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/XOR_2/out addersubtractor_0/fulladder_2/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1101 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/XOR_2/out vdd addersubtractor_0/fulladder_2/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1102 gnd enableblock_0/B_out3 addersubtractor_0/fulladder_2/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1103 vdd enableblock_0/B_out3 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/fulladder_2/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1104 addersubtractor_0/fulladder_2/OR_0/in2 addersubtractor_0/fulladder_2/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1105 addersubtractor_0/fulladder_2/OR_0/in2 addersubtractor_0/fulladder_2/AND_0/not_0/in vdd addersubtractor_0/fulladder_2/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1106 addersubtractor_0/fulladder_2/AND_1/not_0/in addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_2/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1107 addersubtractor_0/fulladder_2/AND_1/not_0/in addersubtractor_0/fulladder_1/C vdd addersubtractor_0/fulladder_2/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1108 gnd addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1109 vdd addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/AND_1/not_0/in addersubtractor_0/fulladder_2/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 addersubtractor_0/fulladder_2/OR_0/in1 addersubtractor_0/fulladder_2/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1111 addersubtractor_0/fulladder_2/OR_0/in1 addersubtractor_0/fulladder_2/AND_1/not_0/in vdd addersubtractor_0/fulladder_2/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1112 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 enableblock_0/B_out3 addersubtractor_0/fulladder_2/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1113 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 enableblock_0/B_out3 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1114 gnd addersubtractor_0/XOR_2/out addersubtractor_0/fulladder_2/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 vdd addersubtractor_0/XOR_2/out addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 enableblock_0/B_out3 addersubtractor_0/fulladder_2/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1117 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 enableblock_0/B_out3 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1118 gnd addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1121 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1122 gnd addersubtractor_0/XOR_2/out addersubtractor_0/fulladder_2/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 vdd addersubtractor_0/XOR_2/out addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1125 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1126 gnd addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1127 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_2/OR_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1129 addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_2/OR_0/NOT_0/in vdd addersubtractor_0/fulladder_2/OR_0/NOT_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1130 addersubtractor_0/fulladder_2/OR_0/NOT_0/in addersubtractor_0/fulladder_2/OR_0/in1 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1131 addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_2/OR_0/in1 vdd addersubtractor_0/fulladder_2/OR_0/NOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1132 gnd addersubtractor_0/fulladder_2/OR_0/in2 addersubtractor_0/fulladder_2/OR_0/NOT_0/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 addersubtractor_0/fulladder_2/OR_0/NOT_0/in addersubtractor_0/fulladder_2/OR_0/in2 addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_2/OR_0/NOR_0/w_32_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1134 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_2/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1135 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/C vdd addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1136 gnd addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1137 vdd addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1138 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_2/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1139 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_1/C vdd addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1140 gnd addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1143 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1144 gnd addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1145 vdd addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 adder2 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1147 adder2 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1148 gnd addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1149 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 adder2 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1150 addersubtractor_0/XOR_0/NAND_2/in1 enableblock_0/A_out2 addersubtractor_0/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1151 addersubtractor_0/XOR_0/NAND_2/in1 enableblock_0/A_out2 vdd addersubtractor_0/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1152 gnd S0 addersubtractor_0/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1153 vdd S0 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1154 addersubtractor_0/XOR_0/NAND_3/in1 enableblock_0/A_out2 addersubtractor_0/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1155 addersubtractor_0/XOR_0/NAND_3/in1 enableblock_0/A_out2 vdd addersubtractor_0/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1156 gnd addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1157 vdd addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_3/in1 addersubtractor_0/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 addersubtractor_0/XOR_0/NAND_3/in2 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1159 addersubtractor_0/XOR_0/NAND_3/in2 addersubtractor_0/XOR_0/NAND_2/in1 vdd addersubtractor_0/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1160 gnd S0 addersubtractor_0/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1161 vdd S0 addersubtractor_0/XOR_0/NAND_3/in2 addersubtractor_0/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 addersubtractor_0/XOR_0/out addersubtractor_0/XOR_0/NAND_3/in1 addersubtractor_0/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1163 addersubtractor_0/XOR_0/out addersubtractor_0/XOR_0/NAND_3/in1 vdd addersubtractor_0/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1164 gnd addersubtractor_0/XOR_0/NAND_3/in2 addersubtractor_0/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 vdd addersubtractor_0/XOR_0/NAND_3/in2 addersubtractor_0/XOR_0/out addersubtractor_0/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 addersubtractor_0/fulladder_3/AND_0/not_0/in addersubtractor_0/XOR_3/out addersubtractor_0/fulladder_3/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1167 addersubtractor_0/fulladder_3/AND_0/not_0/in addersubtractor_0/XOR_3/out vdd addersubtractor_0/fulladder_3/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1168 gnd enableblock_0/B_out1 addersubtractor_0/fulladder_3/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1169 vdd enableblock_0/B_out1 addersubtractor_0/fulladder_3/AND_0/not_0/in addersubtractor_0/fulladder_3/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1171 addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/AND_0/not_0/in vdd addersubtractor_0/fulladder_3/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1172 addersubtractor_0/fulladder_3/AND_1/not_0/in addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_3/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1173 addersubtractor_0/fulladder_3/AND_1/not_0/in addersubtractor_0/fulladder_2/C vdd addersubtractor_0/fulladder_3/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1174 gnd addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 vdd addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/AND_1/not_0/in addersubtractor_0/fulladder_3/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 addersubtractor_0/fulladder_3/OR_0/in1 addersubtractor_0/fulladder_3/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1177 addersubtractor_0/fulladder_3/OR_0/in1 addersubtractor_0/fulladder_3/AND_1/not_0/in vdd addersubtractor_0/fulladder_3/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1178 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 enableblock_0/B_out1 addersubtractor_0/fulladder_3/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1179 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 enableblock_0/B_out1 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1180 gnd addersubtractor_0/XOR_3/out addersubtractor_0/fulladder_3/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1181 vdd addersubtractor_0/XOR_3/out addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1182 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 enableblock_0/B_out1 addersubtractor_0/fulladder_3/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1183 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 enableblock_0/B_out1 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1184 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1185 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1186 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1187 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1188 gnd addersubtractor_0/XOR_3/out addersubtractor_0/fulladder_3/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 vdd addersubtractor_0/XOR_3/out addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1190 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1191 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1192 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1193 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 AND_0/in1 addersubtractor_0/fulladder_3/OR_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1195 AND_0/in1 addersubtractor_0/fulladder_3/OR_0/NOT_0/in vdd addersubtractor_0/fulladder_3/OR_0/NOT_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1196 addersubtractor_0/fulladder_3/OR_0/NOT_0/in addersubtractor_0/fulladder_3/OR_0/in1 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1197 addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_3/OR_0/in1 vdd addersubtractor_0/fulladder_3/OR_0/NOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1198 gnd addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/OR_0/NOT_0/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1199 addersubtractor_0/fulladder_3/OR_0/NOT_0/in addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_3/OR_0/NOR_0/w_32_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1200 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_3/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1201 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/C vdd addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1202 gnd addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1203 vdd addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1204 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_3/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1205 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_2/C vdd addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1206 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1209 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1210 gnd addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1211 vdd addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 adder3 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1213 adder3 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1214 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 adder3 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 addersubtractor_0/XOR_1/NAND_2/in1 enableblock_0/A_out0 addersubtractor_0/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1217 addersubtractor_0/XOR_1/NAND_2/in1 enableblock_0/A_out0 vdd addersubtractor_0/XOR_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1218 gnd S0 addersubtractor_0/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1219 vdd S0 addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1220 addersubtractor_0/XOR_1/NAND_3/in1 enableblock_0/A_out0 addersubtractor_0/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1221 addersubtractor_0/XOR_1/NAND_3/in1 enableblock_0/A_out0 vdd addersubtractor_0/XOR_1/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1222 gnd addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 vdd addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_3/in1 addersubtractor_0/XOR_1/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1224 addersubtractor_0/XOR_1/NAND_3/in2 addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1225 addersubtractor_0/XOR_1/NAND_3/in2 addersubtractor_0/XOR_1/NAND_2/in1 vdd addersubtractor_0/XOR_1/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1226 gnd S0 addersubtractor_0/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 vdd S0 addersubtractor_0/XOR_1/NAND_3/in2 addersubtractor_0/XOR_1/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 addersubtractor_0/XOR_1/out addersubtractor_0/XOR_1/NAND_3/in1 addersubtractor_0/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1229 addersubtractor_0/XOR_1/out addersubtractor_0/XOR_1/NAND_3/in1 vdd addersubtractor_0/XOR_1/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1230 gnd addersubtractor_0/XOR_1/NAND_3/in2 addersubtractor_0/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1231 vdd addersubtractor_0/XOR_1/NAND_3/in2 addersubtractor_0/XOR_1/out addersubtractor_0/XOR_1/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 addersubtractor_0/XOR_2/NAND_2/in1 enableblock_0/B_out2 addersubtractor_0/XOR_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1233 addersubtractor_0/XOR_2/NAND_2/in1 enableblock_0/B_out2 vdd addersubtractor_0/XOR_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1234 gnd S0 addersubtractor_0/XOR_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1235 vdd S0 addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1236 addersubtractor_0/XOR_2/NAND_3/in1 enableblock_0/B_out2 addersubtractor_0/XOR_2/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1237 addersubtractor_0/XOR_2/NAND_3/in1 enableblock_0/B_out2 vdd addersubtractor_0/XOR_2/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1238 gnd addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 vdd addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_3/in1 addersubtractor_0/XOR_2/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1240 addersubtractor_0/XOR_2/NAND_3/in2 addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1241 addersubtractor_0/XOR_2/NAND_3/in2 addersubtractor_0/XOR_2/NAND_2/in1 vdd addersubtractor_0/XOR_2/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1242 gnd S0 addersubtractor_0/XOR_2/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1243 vdd S0 addersubtractor_0/XOR_2/NAND_3/in2 addersubtractor_0/XOR_2/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1244 addersubtractor_0/XOR_2/out addersubtractor_0/XOR_2/NAND_3/in1 addersubtractor_0/XOR_2/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1245 addersubtractor_0/XOR_2/out addersubtractor_0/XOR_2/NAND_3/in1 vdd addersubtractor_0/XOR_2/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1246 gnd addersubtractor_0/XOR_2/NAND_3/in2 addersubtractor_0/XOR_2/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1247 vdd addersubtractor_0/XOR_2/NAND_3/in2 addersubtractor_0/XOR_2/out addersubtractor_0/XOR_2/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1248 addersubtractor_0/XOR_3/NAND_2/in1 enableblock_0/B_out0 addersubtractor_0/XOR_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1249 addersubtractor_0/XOR_3/NAND_2/in1 enableblock_0/B_out0 vdd addersubtractor_0/XOR_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1250 gnd S0 addersubtractor_0/XOR_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 vdd S0 addersubtractor_0/XOR_3/NAND_2/in1 addersubtractor_0/XOR_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1252 addersubtractor_0/XOR_3/NAND_3/in1 enableblock_0/B_out0 addersubtractor_0/XOR_3/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1253 addersubtractor_0/XOR_3/NAND_3/in1 enableblock_0/B_out0 vdd addersubtractor_0/XOR_3/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1254 gnd addersubtractor_0/XOR_3/NAND_2/in1 addersubtractor_0/XOR_3/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1255 vdd addersubtractor_0/XOR_3/NAND_2/in1 addersubtractor_0/XOR_3/NAND_3/in1 addersubtractor_0/XOR_3/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 addersubtractor_0/XOR_3/NAND_3/in2 addersubtractor_0/XOR_3/NAND_2/in1 addersubtractor_0/XOR_3/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1257 addersubtractor_0/XOR_3/NAND_3/in2 addersubtractor_0/XOR_3/NAND_2/in1 vdd addersubtractor_0/XOR_3/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1258 gnd S0 addersubtractor_0/XOR_3/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1259 vdd S0 addersubtractor_0/XOR_3/NAND_3/in2 addersubtractor_0/XOR_3/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1260 addersubtractor_0/XOR_3/out addersubtractor_0/XOR_3/NAND_3/in1 addersubtractor_0/XOR_3/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1261 addersubtractor_0/XOR_3/out addersubtractor_0/XOR_3/NAND_3/in1 vdd addersubtractor_0/XOR_3/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1262 gnd addersubtractor_0/XOR_3/NAND_3/in2 addersubtractor_0/XOR_3/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1263 vdd addersubtractor_0/XOR_3/NAND_3/in2 addersubtractor_0/XOR_3/out addersubtractor_0/XOR_3/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1264 AND_0/not_0/in AND_0/in1 AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1265 AND_0/not_0/in AND_0/in1 vdd AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1266 gnd OR_0/out AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1267 vdd OR_0/out AND_0/not_0/in AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1268 XOR_0/in1 AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1269 XOR_0/in1 AND_0/not_0/in vdd AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1270 AND_1/not_0/in AND_2/in2 AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1271 AND_1/not_0/in AND_2/in2 vdd AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1272 gnd AND_1/in2 AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1273 vdd AND_1/in2 AND_1/not_0/in AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1274 lesser AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1275 lesser AND_1/not_0/in vdd AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1276 AND_2/not_0/in AND_2/in1 AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1277 AND_2/not_0/in AND_2/in1 vdd AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1278 gnd AND_2/in2 AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1279 vdd AND_2/in2 AND_2/not_0/in AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1280 equal AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1281 equal AND_2/not_0/in vdd AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1282 enableblock_1/enable1_1/AND_0/not_0/in A1 enableblock_1/enable1_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1283 enableblock_1/enable1_1/AND_0/not_0/in A1 vdd enableblock_1/enable1_1/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1284 gnd AND_2/in2 enableblock_1/enable1_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1285 vdd AND_2/in2 enableblock_1/enable1_1/AND_0/not_0/in enableblock_1/enable1_1/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1286 comparator_0/A1 enableblock_1/enable1_1/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1287 comparator_0/A1 enableblock_1/enable1_1/AND_0/not_0/in vdd enableblock_1/enable1_1/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1288 enableblock_1/enable1_1/AND_1/not_0/in AND_2/in2 enableblock_1/enable1_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1289 enableblock_1/enable1_1/AND_1/not_0/in AND_2/in2 vdd enableblock_1/enable1_1/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1290 gnd B1 enableblock_1/enable1_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1291 vdd B1 enableblock_1/enable1_1/AND_1/not_0/in enableblock_1/enable1_1/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1292 comparator_0/B1 enableblock_1/enable1_1/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1293 comparator_0/B1 enableblock_1/enable1_1/AND_1/not_0/in vdd enableblock_1/enable1_1/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1294 enableblock_1/enable1_1/AND_2/not_0/in A0 enableblock_1/enable1_1/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1295 enableblock_1/enable1_1/AND_2/not_0/in A0 vdd enableblock_1/enable1_1/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1296 gnd AND_2/in2 enableblock_1/enable1_1/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1297 vdd AND_2/in2 enableblock_1/enable1_1/AND_2/not_0/in enableblock_1/enable1_1/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1298 comparator_0/A0 enableblock_1/enable1_1/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1299 comparator_0/A0 enableblock_1/enable1_1/AND_2/not_0/in vdd enableblock_1/enable1_1/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1300 enableblock_1/enable1_1/AND_3/not_0/in AND_2/in2 enableblock_1/enable1_1/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1301 enableblock_1/enable1_1/AND_3/not_0/in AND_2/in2 vdd enableblock_1/enable1_1/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1302 gnd B0 enableblock_1/enable1_1/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1303 vdd B0 enableblock_1/enable1_1/AND_3/not_0/in enableblock_1/enable1_1/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1304 comparator_0/B0 enableblock_1/enable1_1/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1305 comparator_0/B0 enableblock_1/enable1_1/AND_3/not_0/in vdd enableblock_1/enable1_1/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=45 pd=38 as=0 ps=0
M1306 enableblock_1/enable1_0/AND_0/not_0/in A3 enableblock_1/enable1_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1307 enableblock_1/enable1_0/AND_0/not_0/in A3 vdd enableblock_1/enable1_0/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1308 gnd AND_2/in2 enableblock_1/enable1_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1309 vdd AND_2/in2 enableblock_1/enable1_0/AND_0/not_0/in enableblock_1/enable1_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1310 comparator_0/A3 enableblock_1/enable1_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1311 comparator_0/A3 enableblock_1/enable1_0/AND_0/not_0/in vdd enableblock_1/enable1_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1312 enableblock_1/enable1_0/AND_1/not_0/in AND_2/in2 enableblock_1/enable1_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1313 enableblock_1/enable1_0/AND_1/not_0/in AND_2/in2 vdd enableblock_1/enable1_0/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1314 gnd B3 enableblock_1/enable1_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1315 vdd B3 enableblock_1/enable1_0/AND_1/not_0/in enableblock_1/enable1_0/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1316 comparator_0/B3 enableblock_1/enable1_0/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1317 comparator_0/B3 enableblock_1/enable1_0/AND_1/not_0/in vdd enableblock_1/enable1_0/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1318 enableblock_1/enable1_0/AND_2/not_0/in A2 enableblock_1/enable1_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1319 enableblock_1/enable1_0/AND_2/not_0/in A2 vdd enableblock_1/enable1_0/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1320 gnd AND_2/in2 enableblock_1/enable1_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1321 vdd AND_2/in2 enableblock_1/enable1_0/AND_2/not_0/in enableblock_1/enable1_0/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1322 comparator_0/A2 enableblock_1/enable1_0/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1323 comparator_0/A2 enableblock_1/enable1_0/AND_2/not_0/in vdd enableblock_1/enable1_0/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1324 enableblock_1/enable1_0/AND_3/not_0/in AND_2/in2 enableblock_1/enable1_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1325 enableblock_1/enable1_0/AND_3/not_0/in AND_2/in2 vdd enableblock_1/enable1_0/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1326 gnd B2 enableblock_1/enable1_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1327 vdd B2 enableblock_1/enable1_0/AND_3/not_0/in enableblock_1/enable1_0/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1328 comparator_0/B2 enableblock_1/enable1_0/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1329 comparator_0/B2 enableblock_1/enable1_0/AND_3/not_0/in vdd enableblock_1/enable1_0/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1330 enableblock_0/enable1_1/AND_0/not_0/in A2 enableblock_0/enable1_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1331 enableblock_0/enable1_1/AND_0/not_0/in A2 vdd enableblock_0/enable1_1/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1332 gnd OR_0/out enableblock_0/enable1_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1333 vdd OR_0/out enableblock_0/enable1_1/AND_0/not_0/in enableblock_0/enable1_1/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1334 enableblock_0/B_out3 enableblock_0/enable1_1/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1335 enableblock_0/B_out3 enableblock_0/enable1_1/AND_0/not_0/in vdd enableblock_0/enable1_1/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1336 enableblock_0/enable1_1/AND_1/not_0/in OR_0/out enableblock_0/enable1_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1337 enableblock_0/enable1_1/AND_1/not_0/in OR_0/out vdd enableblock_0/enable1_1/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1338 gnd B2 enableblock_0/enable1_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1339 vdd B2 enableblock_0/enable1_1/AND_1/not_0/in enableblock_0/enable1_1/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1340 enableblock_0/B_out2 enableblock_0/enable1_1/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1341 enableblock_0/B_out2 enableblock_0/enable1_1/AND_1/not_0/in vdd enableblock_0/enable1_1/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1342 enableblock_0/enable1_1/AND_2/not_0/in A3 enableblock_0/enable1_1/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1343 enableblock_0/enable1_1/AND_2/not_0/in A3 vdd enableblock_0/enable1_1/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1344 gnd OR_0/out enableblock_0/enable1_1/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1345 vdd OR_0/out enableblock_0/enable1_1/AND_2/not_0/in enableblock_0/enable1_1/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1346 enableblock_0/B_out1 enableblock_0/enable1_1/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1347 enableblock_0/B_out1 enableblock_0/enable1_1/AND_2/not_0/in vdd enableblock_0/enable1_1/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1348 enableblock_0/enable1_1/AND_3/not_0/in OR_0/out enableblock_0/enable1_1/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1349 enableblock_0/enable1_1/AND_3/not_0/in OR_0/out vdd enableblock_0/enable1_1/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1350 gnd B3 enableblock_0/enable1_1/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1351 vdd B3 enableblock_0/enable1_1/AND_3/not_0/in enableblock_0/enable1_1/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1352 enableblock_0/B_out0 enableblock_0/enable1_1/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1353 enableblock_0/B_out0 enableblock_0/enable1_1/AND_3/not_0/in vdd enableblock_0/enable1_1/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1354 enableblock_0/enable1_0/AND_0/not_0/in A0 enableblock_0/enable1_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1355 enableblock_0/enable1_0/AND_0/not_0/in A0 vdd enableblock_0/enable1_0/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1356 gnd OR_0/out enableblock_0/enable1_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1357 vdd OR_0/out enableblock_0/enable1_0/AND_0/not_0/in enableblock_0/enable1_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1358 enableblock_0/A_out3 enableblock_0/enable1_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1359 enableblock_0/A_out3 enableblock_0/enable1_0/AND_0/not_0/in vdd enableblock_0/enable1_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1360 enableblock_0/enable1_0/AND_1/not_0/in OR_0/out enableblock_0/enable1_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1361 enableblock_0/enable1_0/AND_1/not_0/in OR_0/out vdd enableblock_0/enable1_0/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1362 gnd B0 enableblock_0/enable1_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1363 vdd B0 enableblock_0/enable1_0/AND_1/not_0/in enableblock_0/enable1_0/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1364 enableblock_0/A_out2 enableblock_0/enable1_0/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1365 enableblock_0/A_out2 enableblock_0/enable1_0/AND_1/not_0/in vdd enableblock_0/enable1_0/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1366 enableblock_0/enable1_0/AND_2/not_0/in A1 enableblock_0/enable1_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1367 enableblock_0/enable1_0/AND_2/not_0/in A1 vdd enableblock_0/enable1_0/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1368 gnd OR_0/out enableblock_0/enable1_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1369 vdd OR_0/out enableblock_0/enable1_0/AND_2/not_0/in enableblock_0/enable1_0/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1370 enableblock_0/A_out1 enableblock_0/enable1_0/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1371 enableblock_0/A_out1 enableblock_0/enable1_0/AND_2/not_0/in vdd enableblock_0/enable1_0/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1372 enableblock_0/enable1_0/AND_3/not_0/in OR_0/out enableblock_0/enable1_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1373 enableblock_0/enable1_0/AND_3/not_0/in OR_0/out vdd enableblock_0/enable1_0/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1374 gnd B1 enableblock_0/enable1_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1375 vdd B1 enableblock_0/enable1_0/AND_3/not_0/in enableblock_0/enable1_0/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1376 enableblock_0/A_out0 enableblock_0/enable1_0/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1377 enableblock_0/A_out0 enableblock_0/enable1_0/AND_3/not_0/in vdd enableblock_0/enable1_0/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1378 enableblock_2/enable1_1/AND_0/not_0/in A1 enableblock_2/enable1_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1379 enableblock_2/enable1_1/AND_0/not_0/in A1 vdd enableblock_2/enable1_1/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1380 gnd enableblock_2/En enableblock_2/enable1_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1381 vdd enableblock_2/En enableblock_2/enable1_1/AND_0/not_0/in enableblock_2/enable1_1/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1382 andblock_0/A1 enableblock_2/enable1_1/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1383 andblock_0/A1 enableblock_2/enable1_1/AND_0/not_0/in vdd enableblock_2/enable1_1/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1384 enableblock_2/enable1_1/AND_1/not_0/in enableblock_2/En enableblock_2/enable1_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1385 enableblock_2/enable1_1/AND_1/not_0/in enableblock_2/En vdd enableblock_2/enable1_1/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1386 gnd B1 enableblock_2/enable1_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1387 vdd B1 enableblock_2/enable1_1/AND_1/not_0/in enableblock_2/enable1_1/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1388 andblock_0/B1 enableblock_2/enable1_1/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1389 andblock_0/B1 enableblock_2/enable1_1/AND_1/not_0/in vdd enableblock_2/enable1_1/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1390 enableblock_2/enable1_1/AND_2/not_0/in A0 enableblock_2/enable1_1/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1391 enableblock_2/enable1_1/AND_2/not_0/in A0 vdd enableblock_2/enable1_1/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1392 gnd enableblock_2/En enableblock_2/enable1_1/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1393 vdd enableblock_2/En enableblock_2/enable1_1/AND_2/not_0/in enableblock_2/enable1_1/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1394 andblock_0/A0 enableblock_2/enable1_1/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1395 andblock_0/A0 enableblock_2/enable1_1/AND_2/not_0/in vdd enableblock_2/enable1_1/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1396 enableblock_2/enable1_1/AND_3/not_0/in enableblock_2/En enableblock_2/enable1_1/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1397 enableblock_2/enable1_1/AND_3/not_0/in enableblock_2/En vdd enableblock_2/enable1_1/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1398 gnd B0 enableblock_2/enable1_1/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 vdd B0 enableblock_2/enable1_1/AND_3/not_0/in enableblock_2/enable1_1/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1400 andblock_0/B0 enableblock_2/enable1_1/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1401 andblock_0/B0 enableblock_2/enable1_1/AND_3/not_0/in vdd enableblock_2/enable1_1/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1402 enableblock_2/enable1_0/AND_0/not_0/in A3 enableblock_2/enable1_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1403 enableblock_2/enable1_0/AND_0/not_0/in A3 vdd enableblock_2/enable1_0/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1404 gnd enableblock_2/En enableblock_2/enable1_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1405 vdd enableblock_2/En enableblock_2/enable1_0/AND_0/not_0/in enableblock_2/enable1_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1406 andblock_0/A3 enableblock_2/enable1_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1407 andblock_0/A3 enableblock_2/enable1_0/AND_0/not_0/in vdd enableblock_2/enable1_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1408 enableblock_2/enable1_0/AND_1/not_0/in enableblock_2/En enableblock_2/enable1_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1409 enableblock_2/enable1_0/AND_1/not_0/in enableblock_2/En vdd enableblock_2/enable1_0/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1410 gnd B3 enableblock_2/enable1_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1411 vdd B3 enableblock_2/enable1_0/AND_1/not_0/in enableblock_2/enable1_0/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1412 andblock_0/B3 enableblock_2/enable1_0/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1413 andblock_0/B3 enableblock_2/enable1_0/AND_1/not_0/in vdd enableblock_2/enable1_0/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1414 enableblock_2/enable1_0/AND_2/not_0/in A2 enableblock_2/enable1_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1415 enableblock_2/enable1_0/AND_2/not_0/in A2 vdd enableblock_2/enable1_0/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1416 gnd enableblock_2/En enableblock_2/enable1_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1417 vdd enableblock_2/En enableblock_2/enable1_0/AND_2/not_0/in enableblock_2/enable1_0/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1418 andblock_0/A2 enableblock_2/enable1_0/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1419 andblock_0/A2 enableblock_2/enable1_0/AND_2/not_0/in vdd enableblock_2/enable1_0/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1420 enableblock_2/enable1_0/AND_3/not_0/in enableblock_2/En enableblock_2/enable1_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1421 enableblock_2/enable1_0/AND_3/not_0/in enableblock_2/En vdd enableblock_2/enable1_0/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1422 gnd B2 enableblock_2/enable1_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1423 vdd B2 enableblock_2/enable1_0/AND_3/not_0/in enableblock_2/enable1_0/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1424 andblock_0/B2 enableblock_2/enable1_0/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1425 andblock_0/B2 enableblock_2/enable1_0/AND_3/not_0/in vdd enableblock_2/enable1_0/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1426 twotofourdecoder_0/AND_0/not_0/in S0 twotofourdecoder_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1427 twotofourdecoder_0/AND_0/not_0/in S0 vdd twotofourdecoder_0/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1428 gnd S1 twotofourdecoder_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1429 vdd S1 twotofourdecoder_0/AND_0/not_0/in twotofourdecoder_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1430 enableblock_2/En twotofourdecoder_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1431 enableblock_2/En twotofourdecoder_0/AND_0/not_0/in vdd twotofourdecoder_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1432 twotofourdecoder_0/AND_1/not_0/in S1 twotofourdecoder_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1433 twotofourdecoder_0/AND_1/not_0/in S1 vdd twotofourdecoder_0/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1434 gnd twotofourdecoder_0/not_0/out twotofourdecoder_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1435 vdd twotofourdecoder_0/not_0/out twotofourdecoder_0/AND_1/not_0/in twotofourdecoder_0/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1436 AND_2/in2 twotofourdecoder_0/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1437 AND_2/in2 twotofourdecoder_0/AND_1/not_0/in vdd twotofourdecoder_0/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1438 twotofourdecoder_0/AND_2/not_0/in twotofourdecoder_0/not_0/out twotofourdecoder_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1439 twotofourdecoder_0/AND_2/not_0/in twotofourdecoder_0/not_0/out vdd twotofourdecoder_0/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1440 gnd twotofourdecoder_0/not_1/out twotofourdecoder_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1441 vdd twotofourdecoder_0/not_1/out twotofourdecoder_0/AND_2/not_0/in twotofourdecoder_0/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1442 OR_0/in2 twotofourdecoder_0/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1443 OR_0/in2 twotofourdecoder_0/AND_2/not_0/in vdd twotofourdecoder_0/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1444 twotofourdecoder_0/AND_3/not_0/in twotofourdecoder_0/not_1/out twotofourdecoder_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1445 twotofourdecoder_0/AND_3/not_0/in twotofourdecoder_0/not_1/out vdd twotofourdecoder_0/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1446 gnd S0 twotofourdecoder_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1447 vdd S0 twotofourdecoder_0/AND_3/not_0/in twotofourdecoder_0/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1448 OR_0/in1 twotofourdecoder_0/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1449 OR_0/in1 twotofourdecoder_0/AND_3/not_0/in vdd twotofourdecoder_0/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1450 twotofourdecoder_0/not_0/out S0 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1451 twotofourdecoder_0/not_0/out S0 vdd twotofourdecoder_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1452 twotofourdecoder_0/not_1/out S1 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1453 twotofourdecoder_0/not_1/out S1 vdd twotofourdecoder_0/not_1/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1454 comparator_0/fourinputOR_0/not_0/in comparator_0/fourinputOR_0/in4 gnd Gnd CMOSN w=4 l=2
+  ad=80 pd=72 as=0 ps=0
M1455 comparator_0/fourinputOR_0/not_0/in comparator_0/AND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1456 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# comparator_0/fourinputOR_0/in3 comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_64_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1457 comparator_0/fourinputOR_0/not_0/in comparator_0/fourinputOR_0/in3 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1458 comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# comparator_0/AND_0/out vdd comparator_0/fourinputOR_0/fourinputNOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1459 comparator_0/fourinputOR_0/not_0/in comparator_0/fourinputOR_0/in4 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_97_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1460 gnd comparator_0/fourinputOR_0/in2 comparator_0/fourinputOR_0/not_0/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1461 comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# comparator_0/fourinputOR_0/in2 comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1462 greater comparator_0/fourinputOR_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1463 greater comparator_0/fourinputOR_0/not_0/in vdd comparator_0/fourinputOR_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1464 comparator_0/AND_0/not_0/in comparator_0/not_0/out comparator_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1465 comparator_0/AND_0/not_0/in comparator_0/not_0/out vdd comparator_0/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1466 gnd comparator_0/A3 comparator_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1467 vdd comparator_0/A3 comparator_0/AND_0/not_0/in comparator_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1468 comparator_0/AND_0/out comparator_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1469 comparator_0/AND_0/out comparator_0/AND_0/not_0/in vdd comparator_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1470 comparator_0/not_0/out comparator_0/B3 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1471 comparator_0/not_0/out comparator_0/B3 vdd comparator_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1472 comparator_0/not_1/out comparator_0/B2 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1473 comparator_0/not_1/out comparator_0/B2 vdd comparator_0/not_1/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1474 comparator_0/not_2/out comparator_0/B1 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1475 comparator_0/not_2/out comparator_0/B1 vdd comparator_0/not_2/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1476 comparator_0/not_3/out comparator_0/B0 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1477 comparator_0/not_3/out comparator_0/B0 vdd comparator_0/not_3/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1478 comparator_0/fourinputOR_0/in3 comparator_0/fourinputAND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1479 comparator_0/fourinputOR_0/in3 comparator_0/fourinputAND_0/not_0/in vdd comparator_0/fourinputAND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1480 comparator_0/fourinputAND_0/not_0/in comparator_0/not_2/out comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1481 gnd comparator_0/XNOR_0/out comparator_0/fourinputAND_0/fourinputNAND_0/a_76_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1482 comparator_0/fourinputAND_0/not_0/in comparator_0/XNOR_1/out vdd comparator_0/fourinputAND_0/fourinputNAND_0/w_63_0# CMOSP w=4 l=2
+  ad=80 pd=72 as=0 ps=0
M1483 comparator_0/fourinputAND_0/not_0/in comparator_0/not_2/out vdd comparator_0/fourinputAND_0/fourinputNAND_0/w_0_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1484 comparator_0/fourinputAND_0/fourinputNAND_0/a_76_n14# comparator_0/XNOR_1/out comparator_0/fourinputAND_0/fourinputNAND_0/a_45_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1485 comparator_0/fourinputAND_0/fourinputNAND_0/a_45_n14# comparator_0/A1 comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1486 vdd comparator_0/A1 comparator_0/fourinputAND_0/not_0/in comparator_0/fourinputAND_0/fourinputNAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1487 vdd comparator_0/XNOR_0/out comparator_0/fourinputAND_0/not_0/in comparator_0/fourinputAND_0/fourinputNAND_0/w_100_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1488 AND_2/in1 comparator_0/fourinputAND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1489 AND_2/in1 comparator_0/fourinputAND_1/not_0/in vdd comparator_0/fourinputAND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1490 comparator_0/fourinputAND_1/not_0/in comparator_0/XNOR_3/out comparator_0/fourinputAND_1/fourinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1491 gnd comparator_0/XNOR_2/out comparator_0/fourinputAND_1/fourinputNAND_0/a_76_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1492 comparator_0/fourinputAND_1/not_0/in comparator_0/XNOR_1/out vdd comparator_0/fourinputAND_1/fourinputNAND_0/w_63_0# CMOSP w=4 l=2
+  ad=80 pd=72 as=0 ps=0
M1493 comparator_0/fourinputAND_1/not_0/in comparator_0/XNOR_3/out vdd comparator_0/fourinputAND_1/fourinputNAND_0/w_0_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1494 comparator_0/fourinputAND_1/fourinputNAND_0/a_76_n14# comparator_0/XNOR_1/out comparator_0/fourinputAND_1/fourinputNAND_0/a_45_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1495 comparator_0/fourinputAND_1/fourinputNAND_0/a_45_n14# comparator_0/XNOR_0/out comparator_0/fourinputAND_1/fourinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1496 vdd comparator_0/XNOR_0/out comparator_0/fourinputAND_1/not_0/in comparator_0/fourinputAND_1/fourinputNAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1497 vdd comparator_0/XNOR_2/out comparator_0/fourinputAND_1/not_0/in comparator_0/fourinputAND_1/fourinputNAND_0/w_100_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1498 comparator_0/threeinputAND_0/not_0/in comparator_0/not_1/out comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1499 comparator_0/threeinputAND_0/not_0/in comparator_0/XNOR_0/out vdd comparator_0/threeinputAND_0/threeinputNAND_0/w_63_0# CMOSP w=4 l=2
+  ad=60 pd=54 as=0 ps=0
M1500 comparator_0/threeinputAND_0/not_0/in comparator_0/not_1/out vdd comparator_0/threeinputAND_0/threeinputNAND_0/w_0_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1501 gnd comparator_0/XNOR_0/out comparator_0/threeinputAND_0/threeinputNAND_0/a_45_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1502 comparator_0/threeinputAND_0/threeinputNAND_0/a_45_n14# comparator_0/A2 comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1503 vdd comparator_0/A2 comparator_0/threeinputAND_0/not_0/in comparator_0/threeinputAND_0/threeinputNAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1504 comparator_0/fourinputOR_0/in2 comparator_0/threeinputAND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1505 comparator_0/fourinputOR_0/in2 comparator_0/threeinputAND_0/not_0/in vdd comparator_0/threeinputAND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1506 comparator_0/fourinputOR_0/in4 comparator_0/fiveinputAND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1507 comparator_0/fourinputOR_0/in4 comparator_0/fiveinputAND_0/not_0/in vdd comparator_0/fiveinputAND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1508 comparator_0/fiveinputAND_0/not_0/in comparator_0/not_3/out comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1509 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_113_n14# comparator_0/XNOR_0/out comparator_0/fiveinputAND_0/fiveinputNAND_0/a_76_n14# Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1510 comparator_0/fiveinputAND_0/not_0/in comparator_0/XNOR_2/out vdd comparator_0/fiveinputAND_0/fiveinputNAND_0/w_133_0# CMOSP w=4 l=2
+  ad=100 pd=90 as=0 ps=0
M1511 comparator_0/fiveinputAND_0/not_0/in comparator_0/XNOR_1/out vdd comparator_0/fiveinputAND_0/fiveinputNAND_0/w_63_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1512 comparator_0/fiveinputAND_0/not_0/in comparator_0/not_3/out vdd comparator_0/fiveinputAND_0/fiveinputNAND_0/w_0_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1513 gnd comparator_0/XNOR_2/out comparator_0/fiveinputAND_0/fiveinputNAND_0/a_113_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1514 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_76_n14# comparator_0/XNOR_1/out comparator_0/fiveinputAND_0/fiveinputNAND_0/a_45_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1515 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_45_n14# comparator_0/A0 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1516 vdd comparator_0/A0 comparator_0/fiveinputAND_0/not_0/in comparator_0/fiveinputAND_0/fiveinputNAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1517 vdd comparator_0/XNOR_0/out comparator_0/fiveinputAND_0/not_0/in comparator_0/fiveinputAND_0/fiveinputNAND_0/w_100_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1518 comparator_0/XNOR_1/out comparator_0/XNOR_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1519 comparator_0/XNOR_1/out comparator_0/XNOR_1/not_0/in vdd comparator_0/XNOR_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1520 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/A2 comparator_0/XNOR_1/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1521 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/A2 vdd comparator_0/XNOR_1/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1522 gnd comparator_0/B2 comparator_0/XNOR_1/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1523 vdd comparator_0/B2 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1524 comparator_0/XNOR_1/XOR_0/NAND_3/in1 comparator_0/A2 comparator_0/XNOR_1/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1525 comparator_0/XNOR_1/XOR_0/NAND_3/in1 comparator_0/A2 vdd comparator_0/XNOR_1/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1526 gnd comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1527 vdd comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_3/in1 comparator_0/XNOR_1/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1528 comparator_0/XNOR_1/XOR_0/NAND_3/in2 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1529 comparator_0/XNOR_1/XOR_0/NAND_3/in2 comparator_0/XNOR_1/XOR_0/NAND_2/in1 vdd comparator_0/XNOR_1/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1530 gnd comparator_0/B2 comparator_0/XNOR_1/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1531 vdd comparator_0/B2 comparator_0/XNOR_1/XOR_0/NAND_3/in2 comparator_0/XNOR_1/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1532 comparator_0/XNOR_1/not_0/in comparator_0/XNOR_1/XOR_0/NAND_3/in1 comparator_0/XNOR_1/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1533 comparator_0/XNOR_1/not_0/in comparator_0/XNOR_1/XOR_0/NAND_3/in1 vdd comparator_0/XNOR_1/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1534 gnd comparator_0/XNOR_1/XOR_0/NAND_3/in2 comparator_0/XNOR_1/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1535 vdd comparator_0/XNOR_1/XOR_0/NAND_3/in2 comparator_0/XNOR_1/not_0/in comparator_0/XNOR_1/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1536 comparator_0/XNOR_0/out comparator_0/XNOR_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1537 comparator_0/XNOR_0/out comparator_0/XNOR_0/not_0/in vdd comparator_0/XNOR_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1538 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/A3 comparator_0/XNOR_0/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1539 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/A3 vdd comparator_0/XNOR_0/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1540 gnd comparator_0/B3 comparator_0/XNOR_0/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1541 vdd comparator_0/B3 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1542 comparator_0/XNOR_0/XOR_0/NAND_3/in1 comparator_0/A3 comparator_0/XNOR_0/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1543 comparator_0/XNOR_0/XOR_0/NAND_3/in1 comparator_0/A3 vdd comparator_0/XNOR_0/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1544 gnd comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1545 vdd comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_3/in1 comparator_0/XNOR_0/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1546 comparator_0/XNOR_0/XOR_0/NAND_3/in2 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1547 comparator_0/XNOR_0/XOR_0/NAND_3/in2 comparator_0/XNOR_0/XOR_0/NAND_2/in1 vdd comparator_0/XNOR_0/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1548 gnd comparator_0/B3 comparator_0/XNOR_0/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1549 vdd comparator_0/B3 comparator_0/XNOR_0/XOR_0/NAND_3/in2 comparator_0/XNOR_0/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1550 comparator_0/XNOR_0/not_0/in comparator_0/XNOR_0/XOR_0/NAND_3/in1 comparator_0/XNOR_0/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1551 comparator_0/XNOR_0/not_0/in comparator_0/XNOR_0/XOR_0/NAND_3/in1 vdd comparator_0/XNOR_0/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1552 gnd comparator_0/XNOR_0/XOR_0/NAND_3/in2 comparator_0/XNOR_0/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1553 vdd comparator_0/XNOR_0/XOR_0/NAND_3/in2 comparator_0/XNOR_0/not_0/in comparator_0/XNOR_0/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1554 comparator_0/XNOR_2/out comparator_0/XNOR_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1555 comparator_0/XNOR_2/out comparator_0/XNOR_2/not_0/in vdd comparator_0/XNOR_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1556 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/A1 comparator_0/XNOR_2/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1557 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/A1 vdd comparator_0/XNOR_2/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1558 gnd comparator_0/B1 comparator_0/XNOR_2/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1559 vdd comparator_0/B1 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1560 comparator_0/XNOR_2/XOR_0/NAND_3/in1 comparator_0/A1 comparator_0/XNOR_2/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1561 comparator_0/XNOR_2/XOR_0/NAND_3/in1 comparator_0/A1 vdd comparator_0/XNOR_2/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1562 gnd comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1563 vdd comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_3/in1 comparator_0/XNOR_2/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1564 comparator_0/XNOR_2/XOR_0/NAND_3/in2 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1565 comparator_0/XNOR_2/XOR_0/NAND_3/in2 comparator_0/XNOR_2/XOR_0/NAND_2/in1 vdd comparator_0/XNOR_2/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1566 gnd comparator_0/B1 comparator_0/XNOR_2/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1567 vdd comparator_0/B1 comparator_0/XNOR_2/XOR_0/NAND_3/in2 comparator_0/XNOR_2/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1568 comparator_0/XNOR_2/not_0/in comparator_0/XNOR_2/XOR_0/NAND_3/in1 comparator_0/XNOR_2/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1569 comparator_0/XNOR_2/not_0/in comparator_0/XNOR_2/XOR_0/NAND_3/in1 vdd comparator_0/XNOR_2/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1570 gnd comparator_0/XNOR_2/XOR_0/NAND_3/in2 comparator_0/XNOR_2/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1571 vdd comparator_0/XNOR_2/XOR_0/NAND_3/in2 comparator_0/XNOR_2/not_0/in comparator_0/XNOR_2/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1572 comparator_0/XNOR_3/out comparator_0/XNOR_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1573 comparator_0/XNOR_3/out comparator_0/XNOR_3/not_0/in vdd comparator_0/XNOR_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1574 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/A0 comparator_0/XNOR_3/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1575 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/A0 vdd comparator_0/XNOR_3/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1576 gnd comparator_0/B0 comparator_0/XNOR_3/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1577 vdd comparator_0/B0 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1578 comparator_0/XNOR_3/XOR_0/NAND_3/in1 comparator_0/A0 comparator_0/XNOR_3/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1579 comparator_0/XNOR_3/XOR_0/NAND_3/in1 comparator_0/A0 vdd comparator_0/XNOR_3/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1580 gnd comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1581 vdd comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_3/in1 comparator_0/XNOR_3/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1582 comparator_0/XNOR_3/XOR_0/NAND_3/in2 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1583 comparator_0/XNOR_3/XOR_0/NAND_3/in2 comparator_0/XNOR_3/XOR_0/NAND_2/in1 vdd comparator_0/XNOR_3/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1584 gnd comparator_0/B0 comparator_0/XNOR_3/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1585 vdd comparator_0/B0 comparator_0/XNOR_3/XOR_0/NAND_3/in2 comparator_0/XNOR_3/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1586 comparator_0/XNOR_3/not_0/in comparator_0/XNOR_3/XOR_0/NAND_3/in1 comparator_0/XNOR_3/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1587 comparator_0/XNOR_3/not_0/in comparator_0/XNOR_3/XOR_0/NAND_3/in1 vdd comparator_0/XNOR_3/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1588 gnd comparator_0/XNOR_3/XOR_0/NAND_3/in2 comparator_0/XNOR_3/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1589 vdd comparator_0/XNOR_3/XOR_0/NAND_3/in2 comparator_0/XNOR_3/not_0/in comparator_0/XNOR_3/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1590 AND_1/in2 greater gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1591 comparator_0/NOR_0/a_13_6# greater vdd comparator_0/NOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1592 gnd AND_2/in1 AND_1/in2 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1593 AND_1/in2 AND_2/in1 comparator_0/NOR_0/a_13_6# comparator_0/NOR_0/w_32_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1594 andblock_0/AND_0/not_0/in andblock_0/A3 andblock_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1595 andblock_0/AND_0/not_0/in andblock_0/A3 vdd andblock_0/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1596 gnd andblock_0/B3 andblock_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1597 vdd andblock_0/B3 andblock_0/AND_0/not_0/in andblock_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1598 and3 andblock_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1599 and3 andblock_0/AND_0/not_0/in vdd andblock_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1600 andblock_0/AND_1/not_0/in andblock_0/A2 andblock_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1601 andblock_0/AND_1/not_0/in andblock_0/A2 vdd andblock_0/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1602 gnd andblock_0/B2 andblock_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1603 vdd andblock_0/B2 andblock_0/AND_1/not_0/in andblock_0/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1604 and2 andblock_0/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1605 and2 andblock_0/AND_1/not_0/in vdd andblock_0/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1606 andblock_0/AND_2/not_0/in andblock_0/A1 andblock_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1607 andblock_0/AND_2/not_0/in andblock_0/A1 vdd andblock_0/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1608 gnd andblock_0/B1 andblock_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1609 vdd andblock_0/B1 andblock_0/AND_2/not_0/in andblock_0/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1610 and1 andblock_0/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1611 and1 andblock_0/AND_2/not_0/in vdd andblock_0/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1612 andblock_0/AND_3/not_0/in andblock_0/A0 andblock_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1613 andblock_0/AND_3/not_0/in andblock_0/A0 vdd andblock_0/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1614 gnd andblock_0/B0 andblock_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1615 vdd andblock_0/B0 andblock_0/AND_3/not_0/in andblock_0/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1616 and0 andblock_0/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1617 and0 andblock_0/AND_3/not_0/in vdd andblock_0/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1618 XOR_0/NAND_2/in1 XOR_0/in1 XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1619 XOR_0/NAND_2/in1 XOR_0/in1 vdd XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1620 gnd OR_0/in1 XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1621 vdd OR_0/in1 XOR_0/NAND_2/in1 XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1622 XOR_0/NAND_3/in1 XOR_0/in1 XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1623 XOR_0/NAND_3/in1 XOR_0/in1 vdd XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1624 gnd XOR_0/NAND_2/in1 XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1625 vdd XOR_0/NAND_2/in1 XOR_0/NAND_3/in1 XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1626 XOR_0/NAND_3/in2 XOR_0/NAND_2/in1 XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1627 XOR_0/NAND_3/in2 XOR_0/NAND_2/in1 vdd XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1628 gnd OR_0/in1 XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1629 vdd OR_0/in1 XOR_0/NAND_3/in2 XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1630 Carry XOR_0/NAND_3/in1 XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1631 Carry XOR_0/NAND_3/in1 vdd XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1632 gnd XOR_0/NAND_3/in2 XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1633 vdd XOR_0/NAND_3/in2 Carry XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1634 OR_0/out OR_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1635 OR_0/out OR_0/NOT_0/in vdd OR_0/NOT_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1636 OR_0/NOT_0/in OR_0/in1 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1637 OR_0/NOR_0/a_13_6# OR_0/in1 vdd OR_0/NOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1638 gnd OR_0/in2 OR_0/NOT_0/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1639 OR_0/NOT_0/in OR_0/in2 OR_0/NOR_0/a_13_6# OR_0/NOR_0/w_32_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 comparator_0/A2 comparator_0/XNOR_1/XOR_0/NAND_1/w_0_0# 0.06fF
C1 comparator_0/XNOR_3/out comparator_0/XNOR_3/not_0/w_0_0# 0.03fF
C2 twotofourdecoder_0/AND_0/not_0/in vdd 0.29fF
C3 vdd addersubtractor_0/fulladder_1/AND_0/NAND_0/w_32_0# 0.05fF
C4 OR_0/in2 twotofourdecoder_0/AND_2/not_0/in 0.02fF
C5 addersubtractor_0/fulladder_2/AND_0/not_0/in gnd 0.04fF
C6 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_32_0# 0.06fF
C7 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_32_0# 0.03fF
C8 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_32_0# 0.06fF
C9 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_0_0# 0.03fF
C10 addersubtractor_0/XOR_0/NAND_2/in1 gnd 0.15fF
C11 addersubtractor_0/fulladder_0/OR_0/NOT_0/w_0_0# vdd 0.05fF
C12 twotofourdecoder_0/AND_0/NAND_0/w_32_0# S1 0.06fF
C13 addersubtractor_0/fulladder_2/XOR_0/NAND_0/a_6_n14# gnd 0.57fF
C14 vdd addersubtractor_0/fulladder_2/AND_1/not_0/w_0_0# 0.05fF
C15 vdd addersubtractor_0/fulladder_1/AND_1/not_0/in 0.29fF
C16 twotofourdecoder_0/AND_1/not_0/in vdd 0.29fF
C17 enableblock_0/B_out0 vdd 0.11fF
C18 B2 AND_2/in2 0.06fF
C19 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_1/a_6_n14# 0.57fF
C20 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_32_0# 0.05fF
C21 vdd addersubtractor_0/XOR_0/NAND_1/w_32_0# 0.05fF
C22 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_1/a_6_n14# 0.12fF
C23 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_1/a_6_n14# 0.57fF
C24 enableblock_2/En S0 0.75fF
C25 twotofourdecoder_0/AND_1/not_0/in AND_2/in2 0.02fF
C26 addersubtractor_0/fulladder_3/OR_0/NOT_0/in addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# 0.04fF
C27 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_32_0# 0.05fF
C28 vdd addersubtractor_0/fulladder_1/OR_0/NOR_0/w_0_0# 0.05fF
C29 comparator_0/A3 comparator_0/XNOR_0/XOR_0/NAND_0/w_0_0# 0.06fF
C30 comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# vdd 0.17fF
C31 addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_1/OR_0/NOR_0/w_32_0# 0.03fF
C32 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_0_0# 0.05fF
C33 S1 twotofourdecoder_0/not_0/out 0.14fF
C34 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_1/a_6_n14# 0.12fF
C35 XOR_0/NAND_0/a_6_n14# XOR_0/NAND_2/in1 0.12fF
C36 twotofourdecoder_0/AND_0/not_0/w_0_0# vdd 0.05fF
C37 AND_2/NAND_0/w_0_0# AND_2/not_0/in 0.03fF
C38 enableblock_2/enable1_1/AND_0/not_0/w_0_0# enableblock_2/enable1_1/AND_0/not_0/in 0.06fF
C39 comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# 0.04fF
C40 comparator_0/fourinputOR_0/not_0/w_0_0# comparator_0/fourinputOR_0/not_0/in 0.06fF
C41 comparator_0/A1 comparator_0/XNOR_2/XOR_0/NAND_0/w_0_0# 0.06fF
C42 XOR_0/NAND_3/in1 XOR_0/NAND_1/a_6_n14# 0.12fF
C43 comparator_0/AND_0/not_0/w_0_0# vdd 0.05fF
C44 S1 vdd 0.13fF
C45 enableblock_2/enable1_0/AND_3/NAND_0/w_32_0# enableblock_2/enable1_0/AND_3/not_0/in 0.03fF
C46 andblock_0/B3 andblock_0/AND_0/NAND_0/w_32_0# 0.06fF
C47 gnd addersubtractor_0/XOR_3/NAND_2/in1 0.15fF
C48 vdd addersubtractor_0/XOR_2/NAND_2/w_0_0# 0.05fF
C49 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/fulladder_1/OR_0/in2 0.02fF
C50 addersubtractor_0/XOR_2/out addersubtractor_0/XOR_2/NAND_3/w_0_0# 0.03fF
C51 comparator_0/A0 comparator_0/XNOR_3/XOR_0/NAND_0/w_0_0# 0.06fF
C52 comparator_0/not_0/w_0_0# vdd 0.05fF
C53 enableblock_2/enable1_0/AND_1/NAND_0/w_32_0# vdd 0.05fF
C54 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_63_0# comparator_0/XNOR_1/out 0.06fF
C55 enableblock_2/enable1_1/AND_3/NAND_0/a_6_n14# enableblock_2/enable1_1/AND_3/not_0/in 0.12fF
C56 addersubtractor_0/XOR_1/NAND_3/in1 addersubtractor_0/XOR_1/NAND_3/w_0_0# 0.06fF
C57 enableblock_0/enable1_1/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C58 enableblock_1/enable1_0/AND_3/not_0/w_0_0# vdd 0.05fF
C59 comparator_0/fourinputAND_0/fourinputNAND_0/a_76_n14# comparator_0/XNOR_1/out 0.23fF
C60 enableblock_0/B_out0 addersubtractor_0/XOR_3/NAND_1/w_0_0# 0.06fF
C61 andblock_0/AND_3/not_0/in andblock_0/AND_3/NAND_0/w_32_0# 0.03fF
C62 comparator_0/XNOR_2/not_0/w_0_0# vdd 0.05fF
C63 comparator_0/fourinputAND_1/fourinputNAND_0/w_100_0# comparator_0/fourinputAND_1/not_0/in 0.03fF
C64 comparator_0/XNOR_2/out comparator_0/XNOR_1/out 0.21fF
C65 addersubtractor_0/fulladder_1/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_1/AND_1/not_0/in 0.06fF
C66 XOR_0/NAND_3/in1 vdd 0.25fF
C67 comparator_0/fourinputOR_0/fourinputNOR_0/w_0_0# comparator_0/AND_0/out 0.06fF
C68 enableblock_1/enable1_1/AND_2/NAND_0/a_6_n14# enableblock_1/enable1_1/AND_2/not_0/in 0.12fF
C69 twotofourdecoder_0/AND_1/not_0/w_0_0# twotofourdecoder_0/AND_1/not_0/in 0.06fF
C70 addersubtractor_0/XOR_2/NAND_2/w_0_0# addersubtractor_0/XOR_2/NAND_3/in2 0.03fF
C71 gnd addersubtractor_0/XOR_2/NAND_0/a_6_n14# 0.57fF
C72 comparator_0/XNOR_3/not_0/w_0_0# vdd 0.05fF
C73 twotofourdecoder_0/AND_0/not_0/in twotofourdecoder_0/AND_0/NAND_0/w_0_0# 0.03fF
C74 enableblock_2/enable1_0/AND_0/NAND_0/w_0_0# vdd 0.05fF
C75 comparator_0/fourinputAND_1/not_0/in comparator_0/fourinputAND_1/fourinputNAND_0/a_6_n14# 0.11fF
C76 comparator_0/not_3/w_0_0# comparator_0/not_3/out 0.03fF
C77 enableblock_2/enable1_0/AND_1/NAND_0/a_6_n14# enableblock_2/enable1_0/AND_1/not_0/in 0.12fF
C78 enableblock_0/enable1_1/AND_2/NAND_0/a_6_n14# gnd 0.57fF
C79 enableblock_0/enable1_1/AND_1/not_0/w_0_0# vdd 0.05fF
C80 XOR_0/NAND_1/w_32_0# vdd 0.05fF
C81 comparator_0/NOR_0/w_0_0# vdd 0.05fF
C82 comparator_0/XNOR_1/out gnd 0.69fF
C83 comparator_0/NOR_0/w_32_0# vdd 0.03fF
C84 AND_1/NAND_0/a_6_n14# AND_1/not_0/in 0.12fF
C85 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_0_0# addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 0.03fF
C86 enableblock_0/enable1_1/AND_2/NAND_0/w_0_0# vdd 0.05fF
C87 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_0/w_0_0# 0.03fF
C88 andblock_0/AND_3/not_0/w_0_0# andblock_0/AND_3/not_0/in 0.06fF
C89 enableblock_2/enable1_1/AND_0/not_0/in gnd 0.04fF
C90 S0 addersubtractor_0/XOR_1/NAND_2/w_32_0# 0.06fF
C91 vdd addersubtractor_0/fulladder_1/OR_0/NOT_0/in 0.11fF
C92 twotofourdecoder_0/not_1/out gnd 3.35fF
C93 OR_0/in2 vdd 0.33fF
C94 A0 S0 0.13fF
C95 comparator_0/threeinputAND_0/threeinputNAND_0/w_0_0# comparator_0/not_1/out 0.06fF
C96 enableblock_1/enable1_0/AND_3/NAND_0/a_6_n14# enableblock_1/enable1_0/AND_3/not_0/in 0.12fF
C97 twotofourdecoder_0/AND_3/NAND_0/w_0_0# twotofourdecoder_0/AND_3/not_0/in 0.03fF
C98 andblock_0/B0 andblock_0/AND_3/NAND_0/w_32_0# 0.06fF
C99 andblock_0/B1 andblock_0/AND_2/NAND_0/w_32_0# 0.06fF
C100 addersubtractor_0/fulladder_2/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_2/OR_0/in1 0.03fF
C101 enableblock_1/enable1_0/AND_1/not_0/w_0_0# comparator_0/B3 0.03fF
C102 addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/OR_0/NOT_0/in 0.26fF
C103 vdd addersubtractor_0/XOR_0/NAND_2/w_0_0# 0.05fF
C104 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_0_0# enableblock_0/B_out3 0.06fF
C105 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_32_0# 0.06fF
C106 OR_0/in2 AND_2/in2 1.07fF
C107 twotofourdecoder_0/not_0/w_0_0# S0 0.06fF
C108 enableblock_2/En vdd 0.26fF
C109 enableblock_0/A_out3 S0 0.06fF
C110 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# vdd 0.18fF
C111 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_0_0# 0.05fF
C112 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 0.25fF
C113 addersubtractor_0/fulladder_1/OR_0/NOT_0/in addersubtractor_0/fulladder_1/C 0.02fF
C114 XOR_0/NAND_3/w_0_0# vdd 0.05fF
C115 S0 addersubtractor_0/XOR_3/NAND_2/w_32_0# 0.06fF
C116 comparator_0/AND_0/NAND_0/w_32_0# comparator_0/AND_0/not_0/in 0.03fF
C117 enableblock_2/enable1_0/AND_3/not_0/in gnd 0.04fF
C118 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 0.25fF
C119 vdd addersubtractor_0/fulladder_0/AND_0/not_0/in 0.03fF
C120 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_0/a_6_n14# 0.12fF
C121 andblock_0/A2 enableblock_2/enable1_0/AND_2/not_0/in 0.02fF
C122 OR_0/NOR_0/a_13_6# OR_0/NOT_0/in 0.04fF
C123 comparator_0/fourinputAND_0/fourinputNAND_0/w_32_0# comparator_0/fourinputAND_0/not_0/in 0.03fF
C124 addersubtractor_0/XOR_1/NAND_3/in1 addersubtractor_0/XOR_1/NAND_1/a_6_n14# 0.12fF
C125 B0 S0 0.17fF
C126 enableblock_0/enable1_0/AND_2/NAND_0/w_32_0# vdd 0.05fF
C127 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 gnd 0.15fF
C128 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_0_0# addersubtractor_0/fulladder_1/C 0.06fF
C129 addersubtractor_0/fulladder_0/AND_0/not_0/in vdd 0.29fF
C130 addersubtractor_0/fulladder_3/AND_0/NAND_0/w_32_0# enableblock_0/B_out1 0.06fF
C131 comparator_0/threeinputAND_0/not_0/in comparator_0/threeinputAND_0/threeinputNAND_0/w_32_0# 0.03fF
C132 comparator_0/fourinputAND_1/fourinputNAND_0/w_0_0# comparator_0/fourinputAND_1/not_0/in 0.03fF
C133 equal AND_2/not_0/in 0.02fF
C134 vdd addersubtractor_0/XOR_3/NAND_3/in2 0.25fF
C135 B3 B1 0.19fF
C136 enableblock_0/A_out0 S0 0.06fF
C137 comparator_0/fourinputOR_0/in2 vdd 0.95fF
C138 enableblock_0/enable1_0/AND_2/not_0/in vdd 0.29fF
C139 comparator_0/A1 comparator_0/XNOR_1/out 0.06fF
C140 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_97_0# 0.03fF
C141 comparator_0/A2 vdd 0.20fF
C142 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 0.25fF
C143 comparator_0/A0 comparator_0/XNOR_1/out 0.10fF
C144 comparator_0/XNOR_3/XOR_0/NAND_2/in1 vdd 0.25fF
C145 comparator_0/threeinputAND_0/threeinputNAND_0/w_0_0# vdd 0.05fF
C146 gnd addersubtractor_0/fulladder_3/AND_0/not_0/in 0.04fF
C147 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_32_0# addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 0.06fF
C148 addersubtractor_0/fulladder_0/OR_0/NOT_0/in addersubtractor_0/fulladder_0/OR_0/NOT_0/w_0_0# 0.06fF
C149 comparator_0/XNOR_0/out comparator_0/fiveinputAND_0/fiveinputNAND_0/w_100_0# 0.06fF
C150 comparator_0/XNOR_0/out comparator_0/XNOR_0/not_0/in 0.02fF
C151 comparator_0/fourinputAND_0/fourinputNAND_0/w_0_0# vdd 0.05fF
C152 addersubtractor_0/fulladder_3/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_3/AND_1/not_0/in 0.12fF
C153 B2 A3 0.82fF
C154 enableblock_0/enable1_1/AND_1/NAND_0/w_32_0# vdd 0.05fF
C155 comparator_0/threeinputAND_0/threeinputNAND_0/w_63_0# vdd 0.05fF
C156 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 0.06fF
C157 adder0 addersubtractor_0/fulladder_0/XOR_1/NAND_3/a_6_n14# 0.12fF
C158 comparator_0/fourinputAND_0/fourinputNAND_0/a_76_n14# gnd 0.04fF
C159 enableblock_2/enable1_1/AND_3/NAND_0/w_32_0# vdd 0.05fF
C160 addersubtractor_0/fulladder_3/AND_0/NAND_0/a_6_n14# addersubtractor_0/XOR_3/out 0.07fF
C161 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# comparator_0/fiveinputAND_0/fiveinputNAND_0/a_45_n14# 0.04fF
C162 comparator_0/XNOR_2/out gnd 0.31fF
C163 gnd enableblock_1/enable1_0/AND_1/NAND_0/a_6_n14# 0.57fF
C164 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_133_0# vdd 0.05fF
C165 vdd enableblock_1/enable1_1/AND_2/NAND_0/w_32_0# 0.05fF
C166 addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_3/a_6_n14# 0.12fF
C167 vdd addersubtractor_0/XOR_1/NAND_1/w_32_0# 0.05fF
C168 enableblock_2/enable1_1/AND_3/not_0/in vdd 0.29fF
C169 comparator_0/B3 vdd 0.26fF
C170 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_32_0# adder1 0.03fF
C171 twotofourdecoder_0/AND_1/NAND_0/w_0_0# vdd 0.05fF
C172 comparator_0/fourinputOR_0/fourinputNOR_0/w_64_0# comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# 0.03fF
C173 enableblock_1/enable1_1/AND_2/NAND_0/w_32_0# AND_2/in2 0.06fF
C174 comparator_0/fiveinputAND_0/not_0/in vdd 2.81fF
C175 twotofourdecoder_0/not_0/out twotofourdecoder_0/not_0/w_0_0# 0.03fF
C176 vdd enableblock_1/enable1_1/AND_2/not_0/in 0.29fF
C177 andblock_0/B3 gnd 0.44fF
C178 comparator_0/B1 vdd 0.35fF
C179 twotofourdecoder_0/AND_3/not_0/w_0_0# vdd 0.05fF
C180 enableblock_2/enable1_0/AND_1/not_0/w_0_0# enableblock_2/enable1_0/AND_1/not_0/in 0.06fF
C181 vdd addersubtractor_0/XOR_1/NAND_2/w_32_0# 0.05fF
C182 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_0_0# 0.06fF
C183 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_1/XOR_1/in2 0.03fF
C184 addersubtractor_0/fulladder_0/AND_1/not_0/in gnd 0.04fF
C185 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_0/w_32_0# 0.03fF
C186 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_32_0# 0.05fF
C187 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_2/a_6_n14# 0.59fF
C188 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_0_0# 0.06fF
C189 comparator_0/not_2/w_0_0# vdd 0.05fF
C190 enableblock_1/enable1_0/AND_1/not_0/in enableblock_1/enable1_0/AND_1/NAND_0/w_32_0# 0.03fF
C191 comparator_0/B0 vdd 0.17fF
C192 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_32_0# 0.05fF
C193 S0 addersubtractor_0/XOR_0/NAND_0/w_32_0# 0.06fF
C194 vdd adder1 0.25fF
C195 A3 S1 0.06fF
C196 and1 andblock_0/AND_2/not_0/w_0_0# 0.03fF
C197 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_32_0# 0.05fF
C198 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_2/a_6_n14# 0.59fF
C199 addersubtractor_0/fulladder_0/OR_0/NOR_0/w_32_0# vdd 0.03fF
C200 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_0_0# 0.06fF
C201 vdd addersubtractor_0/fulladder_1/XOR_1/in2 0.47fF
C202 twotofourdecoder_0/not_0/w_0_0# vdd 0.05fF
C203 A0 AND_2/in2 0.06fF
C204 enableblock_0/A_out3 vdd 0.43fF
C205 addersubtractor_0/fulladder_3/AND_1/not_0/in addersubtractor_0/fulladder_3/OR_0/in1 0.02fF
C206 OR_0/out gnd 3.60fF
C207 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_0_0# vdd 0.05fF
C208 OR_0/NOR_0/w_0_0# vdd 0.05fF
C209 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_2/w_0_0# 0.06fF
C210 AND_2/in1 gnd 0.68fF
C211 gnd addersubtractor_0/XOR_3/NAND_2/a_6_n14# 0.59fF
C212 gnd addersubtractor_0/XOR_0/NAND_1/a_6_n14# 0.57fF
C213 comparator_0/XNOR_0/not_0/w_0_0# vdd 0.05fF
C214 vdd addersubtractor_0/XOR_3/NAND_2/w_32_0# 0.05fF
C215 addersubtractor_0/fulladder_3/OR_0/NOR_0/w_0_0# addersubtractor_0/fulladder_3/OR_0/in1 0.06fF
C216 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 gnd 0.15fF
C217 comparator_0/threeinputAND_0/threeinputNAND_0/a_45_n14# gnd 0.04fF
C218 greater vdd 0.39fF
C219 A2 enableblock_2/enable1_0/AND_2/NAND_0/w_0_0# 0.06fF
C220 S1 twotofourdecoder_0/not_1/w_0_0# 0.06fF
C221 enableblock_2/enable1_1/AND_2/NAND_0/w_32_0# enableblock_2/enable1_1/AND_2/not_0/in 0.03fF
C222 vdd AND_1/not_0/in 0.29fF
C223 comparator_0/fourinputOR_0/in3 vdd 0.18fF
C224 vdd addersubtractor_0/fulladder_3/AND_0/NAND_0/w_0_0# 0.05fF
C225 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_0_0# addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 0.03fF
C226 greater AND_2/in2 0.06fF
C227 enableblock_2/enable1_0/AND_3/NAND_0/w_0_0# enableblock_2/enable1_0/AND_3/not_0/in 0.03fF
C228 comparator_0/fourinputOR_0/fourinputNOR_0/w_0_0# vdd 0.05fF
C229 enableblock_0/A_out0 vdd 0.17fF
C230 vdd addersubtractor_0/XOR_2/NAND_3/w_0_0# 0.05fF
C231 comparator_0/XNOR_2/out comparator_0/A1 0.11fF
C232 enableblock_1/enable1_0/AND_2/not_0/in gnd 0.04fF
C233 enableblock_1/enable1_1/AND_1/NAND_0/w_32_0# enableblock_1/enable1_1/AND_1/not_0/in 0.03fF
C234 A3 enableblock_2/enable1_0/AND_0/NAND_0/w_0_0# 0.06fF
C235 comparator_0/A3 gnd 1.24fF
C236 comparator_0/XNOR_2/out comparator_0/A0 0.06fF
C237 vdd addersubtractor_0/XOR_3/NAND_3/in1 0.25fF
C238 andblock_0/A1 andblock_0/AND_2/NAND_0/w_0_0# 0.06fF
C239 enableblock_0/enable1_0/AND_0/NAND_0/a_6_n14# enableblock_0/enable1_0/AND_0/not_0/in 0.12fF
C240 comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_0_0# 0.03fF
C241 andblock_0/A2 andblock_0/AND_1/NAND_0/a_6_n14# 0.02fF
C242 comparator_0/A1 gnd 1.67fF
C243 enableblock_1/enable1_0/AND_0/NAND_0/w_32_0# enableblock_1/enable1_0/AND_0/not_0/in 0.03fF
C244 addersubtractor_0/fulladder_0/XOR_1/NAND_2/a_6_n14# addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 0.12fF
C245 comparator_0/XNOR_0/XOR_0/NAND_0/w_0_0# vdd 0.05fF
C246 vdd addersubtractor_0/fulladder_3/AND_1/NAND_0/w_32_0# 0.05fF
C247 andblock_0/B1 vdd 0.20fF
C248 enableblock_0/enable1_1/AND_2/NAND_0/w_0_0# A3 0.06fF
C249 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_0_0# S0 0.06fF
C250 andblock_0/A3 andblock_0/AND_0/NAND_0/a_6_n14# 0.07fF
C251 comparator_0/A0 gnd 1.10fF
C252 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_0/w_32_0# 0.03fF
C253 enableblock_0/A_out0 enableblock_0/enable1_0/AND_3/not_0/in 0.02fF
C254 comparator_0/XNOR_2/XOR_0/NAND_0/w_0_0# vdd 0.05fF
C255 addersubtractor_0/fulladder_0/XOR_0/NAND_2/a_6_n14# addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 0.12fF
C256 vdd addersubtractor_0/fulladder_1/AND_0/NAND_0/w_0_0# 0.05fF
C257 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_32_0# addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 0.03fF
C258 addersubtractor_0/fulladder_1/OR_0/in2 addersubtractor_0/fulladder_1/OR_0/NOR_0/w_32_0# 0.06fF
C259 enableblock_1/enable1_0/AND_2/NAND_0/w_32_0# enableblock_1/enable1_0/AND_2/not_0/in 0.03fF
C260 comparator_0/XNOR_3/XOR_0/NAND_0/w_0_0# vdd 0.05fF
C261 twotofourdecoder_0/AND_2/NAND_0/w_32_0# twotofourdecoder_0/not_1/out 0.06fF
C262 enableblock_1/enable1_0/AND_3/not_0/w_0_0# comparator_0/B2 0.03fF
C263 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_0/a_6_n14# 0.12fF
C264 A3 enableblock_2/En 0.13fF
C265 addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# vdd 0.21fF
C266 addersubtractor_0/fulladder_0/OR_0/in1 gnd 0.30fF
C267 addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_32_0# addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 0.03fF
C268 addersubtractor_0/fulladder_0/AND_1/not_0/in addersubtractor_0/fulladder_0/OR_0/in1 0.02fF
C269 comparator_0/NOR_0/a_13_6# vdd 0.21fF
C270 enableblock_0/enable1_1/AND_3/not_0/in gnd 0.04fF
C271 comparator_0/B0 enableblock_1/enable1_1/AND_3/not_0/in 0.02fF
C272 comparator_0/fourinputOR_0/fourinputNOR_0/w_64_0# comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# 0.03fF
C273 A2 B2 0.23fF
C274 vdd addersubtractor_0/fulladder_2/AND_0/not_0/in 0.29fF
C275 twotofourdecoder_0/not_1/out S0 0.13fF
C276 S0 addersubtractor_0/XOR_2/NAND_0/w_32_0# 0.06fF
C277 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_32_0# 0.05fF
C278 vdd addersubtractor_0/XOR_0/NAND_2/in1 0.25fF
C279 B0 enableblock_1/enable1_1/AND_3/NAND_0/w_32_0# 0.06fF
C280 B1 enableblock_1/enable1_1/AND_1/NAND_0/w_32_0# 0.06fF
C281 addersubtractor_0/XOR_2/out gnd 0.56fF
C282 twotofourdecoder_0/AND_1/NAND_0/a_6_n14# twotofourdecoder_0/AND_1/not_0/in 0.12fF
C283 addersubtractor_0/XOR_3/NAND_3/in1 addersubtractor_0/XOR_3/NAND_1/w_0_0# 0.03fF
C284 vdd addersubtractor_0/XOR_0/NAND_0/w_32_0# 0.05fF
C285 comparator_0/AND_0/out comparator_0/XNOR_2/out 0.13fF
C286 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_32_0# 0.03fF
C287 twotofourdecoder_0/AND_3/not_0/in OR_0/in1 0.02fF
C288 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_32_0# 0.06fF
C289 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_0_0# 0.03fF
C290 andblock_0/AND_2/not_0/in gnd 0.04fF
C291 addersubtractor_0/fulladder_3/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_2/C 0.06fF
C292 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_32_0# 0.06fF
C293 vdd addersubtractor_0/fulladder_2/OR_0/NOT_0/w_0_0# 0.05fF
C294 enableblock_0/enable1_0/AND_2/NAND_0/a_6_n14# gnd 0.57fF
C295 enableblock_0/enable1_0/AND_1/not_0/w_0_0# vdd 0.05fF
C296 andblock_0/B1 enableblock_2/enable1_1/AND_1/not_0/in 0.02fF
C297 comparator_0/AND_0/out gnd 0.54fF
C298 enableblock_2/enable1_0/AND_3/not_0/w_0_0# andblock_0/B2 0.03fF
C299 addersubtractor_0/fulladder_0/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_0/AND_0/not_0/in 0.06fF
C300 enableblock_0/enable1_1/AND_1/NAND_0/a_6_n14# enableblock_0/enable1_1/AND_1/not_0/in 0.12fF
C301 AND_0/in1 AND_0/NAND_0/w_0_0# 0.06fF
C302 addersubtractor_0/fulladder_3/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_3/OR_0/in2 0.03fF
C303 enableblock_0/enable1_0/AND_2/NAND_0/w_0_0# vdd 0.05fF
C304 addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_2/OR_0/NOR_0/w_32_0# 0.03fF
C305 enableblock_0/enable1_0/AND_1/NAND_0/w_0_0# enableblock_0/enable1_0/AND_1/not_0/in 0.03fF
C306 andblock_0/AND_0/NAND_0/w_32_0# vdd 0.05fF
C307 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_2/C 0.06fF
C308 A2 S1 0.06fF
C309 enableblock_2/enable1_0/AND_1/NAND_0/w_32_0# enableblock_2/enable1_0/AND_1/not_0/in 0.03fF
C310 vdd addersubtractor_0/XOR_3/NAND_2/in1 0.25fF
C311 enableblock_0/enable1_0/AND_2/not_0/w_0_0# enableblock_0/enable1_0/AND_2/not_0/in 0.06fF
C312 addersubtractor_0/XOR_0/NAND_2/w_0_0# addersubtractor_0/XOR_0/NAND_3/in2 0.03fF
C313 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/fulladder_1/AND_0/NAND_0/w_32_0# 0.03fF
C314 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_32_0# addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 0.03fF
C315 enableblock_2/enable1_1/AND_1/NAND_0/w_0_0# enableblock_2/En 0.06fF
C316 A1 enableblock_2/enable1_1/AND_0/NAND_0/a_6_n14# 0.07fF
C317 enableblock_0/enable1_1/AND_0/NAND_0/a_6_n14# enableblock_0/enable1_1/AND_0/not_0/in 0.12fF
C318 gnd AND_1/NAND_0/a_6_n14# 0.57fF
C319 addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_0/OR_0/NOR_0/w_0_0# 0.03fF
C320 enableblock_2/enable1_1/AND_3/NAND_0/a_6_n14# gnd 0.57fF
C321 enableblock_2/enable1_1/AND_2/not_0/w_0_0# vdd 0.05fF
C322 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/fulladder_2/OR_0/in2 0.02fF
C323 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_76_n14# comparator_0/XNOR_1/out 0.12fF
C324 enableblock_0/B_out2 gnd 0.82fF
C325 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 gnd 0.11fF
C326 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_0_0# 0.05fF
C327 gnd enableblock_1/enable1_1/AND_2/NAND_0/a_6_n14# 0.57fF
C328 vdd enableblock_1/enable1_1/AND_1/not_0/w_0_0# 0.05fF
C329 addersubtractor_0/fulladder_0/OR_0/NOT_0/in addersubtractor_0/fulladder_0/OR_0/NOR_0/w_32_0# 0.03fF
C330 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 gnd 0.11fF
C331 enableblock_0/enable1_1/AND_3/NAND_0/w_32_0# enableblock_0/enable1_1/AND_3/not_0/in 0.03fF
C332 A3 A0 0.19fF
C333 enableblock_2/enable1_1/AND_3/NAND_0/w_0_0# vdd 0.05fF
C334 comparator_0/A2 comparator_0/B2 2.42fF
C335 enableblock_0/A_out1 addersubtractor_0/XOR_1/out 0.11fF
C336 addersubtractor_0/fulladder_1/XOR_1/NAND_1/a_6_n14# gnd 0.57fF
C337 comparator_0/XNOR_1/out vdd 0.36fF
C338 addersubtractor_0/fulladder_2/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_2/AND_1/not_0/in 0.06fF
C339 addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_0_0# 0.06fF
C340 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_32_0# 0.05fF
C341 comparator_0/threeinputAND_0/threeinputNAND_0/w_32_0# comparator_0/A2 0.06fF
C342 vdd enableblock_1/enable1_1/AND_2/NAND_0/w_0_0# 0.05fF
C343 addersubtractor_0/fulladder_1/XOR_0/NAND_1/a_6_n14# gnd 0.57fF
C344 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_0_0# addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 0.03fF
C345 twotofourdecoder_0/AND_2/not_0/in gnd 0.04fF
C346 addersubtractor_0/XOR_2/NAND_3/in1 addersubtractor_0/XOR_2/NAND_3/w_0_0# 0.06fF
C347 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_32_0# 0.05fF
C348 and0 andblock_0/AND_3/not_0/w_0_0# 0.03fF
C349 twotofourdecoder_0/AND_3/NAND_0/a_6_n14# twotofourdecoder_0/AND_3/not_0/in 0.12fF
C350 enableblock_2/enable1_1/AND_0/not_0/in vdd 0.29fF
C351 gnd S0 1.94fF
C352 B2 A1 0.19fF
C353 A3 B0 0.19fF
C354 twotofourdecoder_0/not_1/out vdd 0.64fF
C355 vdd addersubtractor_0/XOR_2/NAND_0/w_32_0# 0.05fF
C356 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_3/a_6_n14# 0.57fF
C357 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_32_0# 0.05fF
C358 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_3/a_6_n14# 0.57fF
C359 enableblock_2/enable1_0/AND_3/NAND_0/w_32_0# vdd 0.05fF
C360 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_32_0# 0.05fF
C361 comparator_0/XNOR_1/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_1/not_0/in 0.03fF
C362 comparator_0/fourinputOR_0/fourinputNOR_0/w_64_0# comparator_0/fourinputOR_0/in3 0.06fF
C363 OR_0/out S0 1.74fF
C364 A2 enableblock_2/En 0.13fF
C365 enableblock_1/enable1_0/AND_3/NAND_0/w_32_0# B2 0.06fF
C366 comparator_0/XNOR_3/out gnd 0.10fF
C367 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_0_0# vdd 0.05fF
C368 Carry vdd 0.25fF
C369 enableblock_0/enable1_0/AND_1/not_0/w_0_0# enableblock_0/A_out2 0.03fF
C370 vdd addersubtractor_0/XOR_3/NAND_3/w_32_0# 0.05fF
C371 gnd addersubtractor_0/XOR_3/NAND_3/a_6_n14# 0.57fF
C372 enableblock_2/enable1_0/AND_3/not_0/in vdd 0.29fF
C373 gnd addersubtractor_0/XOR_1/NAND_2/a_6_n14# 0.59fF
C374 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_32_0# comparator_0/fiveinputAND_0/not_0/in 0.03fF
C375 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_32_0# 0.06fF
C376 enableblock_2/enable1_1/AND_0/not_0/w_0_0# vdd 0.05fF
C377 enableblock_2/enable1_1/AND_2/NAND_0/w_0_0# enableblock_2/enable1_1/AND_2/not_0/in 0.03fF
C378 comparator_0/XNOR_0/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_0/not_0/in 0.03fF
C379 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 vdd 0.25fF
C380 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_1/C 0.06fF
C381 addersubtractor_0/XOR_1/out addersubtractor_0/XOR_1/NAND_3/w_32_0# 0.03fF
C382 comparator_0/XNOR_1/XOR_0/NAND_2/in1 gnd 0.15fF
C383 enableblock_2/enable1_1/AND_3/not_0/w_0_0# enableblock_2/enable1_1/AND_3/not_0/in 0.06fF
C384 A1 S1 0.06fF
C385 comparator_0/not_1/out gnd 0.08fF
C386 enableblock_0/enable1_0/AND_0/not_0/w_0_0# enableblock_0/enable1_0/AND_0/not_0/in 0.06fF
C387 enableblock_1/enable1_1/AND_1/NAND_0/w_0_0# enableblock_1/enable1_1/AND_1/not_0/in 0.03fF
C388 OR_0/NOT_0/w_0_0# OR_0/NOT_0/in 0.06fF
C389 gnd addersubtractor_0/XOR_2/NAND_1/a_6_n14# 0.57fF
C390 addersubtractor_0/fulladder_0/OR_0/NOT_0/in addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# 0.04fF
C391 comparator_0/XNOR_0/XOR_0/NAND_0/a_6_n14# gnd 0.57fF
C392 vdd addersubtractor_0/XOR_0/NAND_3/w_0_0# 0.05fF
C393 comparator_0/XNOR_1/XOR_0/NAND_0/w_0_0# comparator_0/A2 0.06fF
C394 XOR_0/NAND_2/in1 XOR_0/NAND_0/w_32_0# 0.03fF
C395 comparator_0/XNOR_2/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_2/not_0/in 0.03fF
C396 comparator_0/AND_0/not_0/w_0_0# comparator_0/AND_0/not_0/in 0.06fF
C397 addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_0/a_6_n14# 0.12fF
C398 addersubtractor_0/XOR_0/out addersubtractor_0/XOR_0/NAND_3/w_32_0# 0.03fF
C399 enableblock_1/enable1_1/AND_2/not_0/w_0_0# enableblock_1/enable1_1/AND_2/not_0/in 0.06fF
C400 enableblock_0/enable1_0/AND_1/NAND_0/w_32_0# vdd 0.05fF
C401 comparator_0/XNOR_2/XOR_0/NAND_0/a_6_n14# gnd 0.57fF
C402 andblock_0/AND_2/not_0/in andblock_0/AND_2/NAND_0/w_32_0# 0.03fF
C403 comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# gnd 0.47fF
C404 vdd addersubtractor_0/fulladder_3/AND_0/not_0/in 0.29fF
C405 andblock_0/AND_0/not_0/w_0_0# vdd 0.05fF
C406 comparator_0/not_3/out comparator_0/B0 0.02fF
C407 enableblock_0/A_out1 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_0_0# 0.06fF
C408 XOR_0/NAND_1/a_6_n14# gnd 0.57fF
C409 comparator_0/XNOR_3/XOR_0/NAND_0/a_6_n14# gnd 0.57fF
C410 comparator_0/fiveinputAND_0/not_0/in comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# 0.11fF
C411 comparator_0/XNOR_3/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_3/not_0/in 0.03fF
C412 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_63_0# vdd 0.05fF
C413 AND_1/NAND_0/w_0_0# AND_1/not_0/in 0.03fF
C414 comparator_0/XNOR_0/out comparator_0/fiveinputAND_0/fiveinputNAND_0/a_113_n14# 0.14fF
C415 XOR_0/in1 AND_0/not_0/w_0_0# 0.03fF
C416 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_32_0# addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 0.06fF
C417 addersubtractor_0/fulladder_1/OR_0/NOT_0/in addersubtractor_0/fulladder_1/OR_0/NOT_0/w_0_0# 0.06fF
C418 twotofourdecoder_0/not_0/out gnd 0.42fF
C419 addersubtractor_0/XOR_0/NAND_2/a_6_n14# addersubtractor_0/XOR_0/NAND_3/in2 0.12fF
C420 XOR_0/NAND_2/in1 XOR_0/NAND_2/w_0_0# 0.06fF
C421 enableblock_0/enable1_0/AND_0/NAND_0/w_0_0# vdd 0.05fF
C422 enableblock_1/enable1_0/AND_2/NAND_0/w_0_0# enableblock_1/enable1_0/AND_2/not_0/in 0.03fF
C423 enableblock_2/enable1_1/AND_0/NAND_0/w_32_0# enableblock_2/En 0.06fF
C424 enableblock_0/enable1_1/AND_2/not_0/in enableblock_0/B_out1 0.02fF
C425 comparator_0/XNOR_2/out vdd 0.48fF
C426 addersubtractor_0/fulladder_0/XOR_1/NAND_0/a_6_n14# gnd 0.57fF
C427 addersubtractor_0/XOR_1/NAND_3/in1 addersubtractor_0/XOR_1/NAND_1/w_0_0# 0.03fF
C428 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_0/a_6_n14# 0.57fF
C429 vdd addersubtractor_0/fulladder_3/AND_1/not_0/w_0_0# 0.05fF
C430 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 0.06fF
C431 OR_0/NOR_0/a_13_6# OR_0/NOR_0/w_0_0# 0.03fF
C432 enableblock_2/enable1_0/AND_0/NAND_0/w_32_0# vdd 0.05fF
C433 enableblock_1/enable1_0/AND_3/not_0/w_0_0# enableblock_1/enable1_0/AND_3/not_0/in 0.06fF
C434 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_32_0# 0.06fF
C435 adder1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/a_6_n14# 0.12fF
C436 addersubtractor_0/XOR_1/NAND_3/w_32_0# addersubtractor_0/XOR_1/NAND_3/in2 0.06fF
C437 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 0.25fF
C438 enableblock_2/enable1_0/AND_0/NAND_0/w_0_0# enableblock_2/enable1_0/AND_0/not_0/in 0.03fF
C439 enableblock_1/enable1_1/AND_0/NAND_0/w_32_0# vdd 0.05fF
C440 vdd gnd 7.31fF
C441 andblock_0/B3 vdd 0.26fF
C442 enableblock_0/enable1_1/AND_3/NAND_0/w_0_0# OR_0/out 0.06fF
C443 enableblock_0/enable1_1/AND_0/not_0/in gnd 0.04fF
C444 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 0.25fF
C445 comparator_0/XNOR_1/XOR_0/NAND_2/w_32_0# comparator_0/XNOR_1/XOR_0/NAND_3/in2 0.03fF
C446 addersubtractor_0/XOR_3/out addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_32_0# 0.06fF
C447 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_0_0# 0.05fF
C448 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_3/a_6_n14# 0.12fF
C449 addersubtractor_0/fulladder_0/AND_1/not_0/in vdd 0.29fF
C450 vdd AND_1/not_0/w_0_0# 0.05fF
C451 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_32_0# adder2 0.03fF
C452 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_32_0# vdd 0.05fF
C453 enableblock_1/enable1_1/AND_0/NAND_0/w_32_0# AND_2/in2 0.06fF
C454 gnd AND_2/in2 3.67fF
C455 A2 A0 0.19fF
C456 gnd AND_2/NAND_0/a_6_n14# 0.57fF
C457 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_0/AND_1/not_0/in 0.03fF
C458 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_0/w_32_0# 0.03fF
C459 addersubtractor_0/fulladder_1/C gnd 1.14fF
C460 enableblock_2/enable1_1/AND_2/not_0/w_0_0# andblock_0/A0 0.03fF
C461 OR_0/out vdd 0.13fF
C462 enableblock_0/A_out0 addersubtractor_0/XOR_1/NAND_0/w_0_0# 0.06fF
C463 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_2/XOR_1/in2 0.03fF
C464 comparator_0/XNOR_0/XOR_0/NAND_2/w_32_0# comparator_0/XNOR_0/XOR_0/NAND_3/in2 0.03fF
C465 A1 enableblock_2/En 0.13fF
C466 AND_2/in1 vdd 0.12fF
C467 enableblock_2/enable1_0/AND_3/NAND_0/a_6_n14# enableblock_2/enable1_0/AND_3/not_0/in 0.12fF
C468 addersubtractor_0/fulladder_3/AND_0/NAND_0/w_0_0# addersubtractor_0/XOR_3/out 0.06fF
C469 comparator_0/XNOR_0/XOR_0/NAND_0/w_32_0# comparator_0/B3 0.06fF
C470 enableblock_0/enable1_0/AND_3/not_0/in gnd 0.04fF
C471 vdd addersubtractor_0/fulladder_2/OR_0/NOR_0/w_32_0# 0.03fF
C472 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 0.25fF
C473 AND_2/in1 AND_2/in2 0.06fF
C474 A2 B0 0.19fF
C475 AND_2/in1 AND_2/NAND_0/a_6_n14# 0.08fF
C476 enableblock_1/enable1_0/AND_2/NAND_0/w_32_0# vdd 0.05fF
C477 enableblock_0/enable1_1/AND_1/not_0/w_0_0# enableblock_0/enable1_1/AND_1/not_0/in 0.06fF
C478 comparator_0/XNOR_2/XOR_0/NAND_2/w_32_0# comparator_0/XNOR_2/XOR_0/NAND_3/in2 0.03fF
C479 comparator_0/fourinputOR_0/fourinputNOR_0/w_32_0# vdd 0.03fF
C480 enableblock_1/enable1_0/AND_2/NAND_0/w_32_0# AND_2/in2 0.06fF
C481 andblock_0/AND_1/NAND_0/w_32_0# vdd 0.05fF
C482 enableblock_1/enable1_0/AND_2/not_0/in vdd 0.29fF
C483 comparator_0/XNOR_2/XOR_0/NAND_0/w_32_0# comparator_0/B1 0.06fF
C484 addersubtractor_0/fulladder_1/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C485 comparator_0/A3 vdd 0.32fF
C486 enableblock_2/enable1_1/AND_1/not_0/in gnd 0.04fF
C487 addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_0_0# addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 0.03fF
C488 comparator_0/XNOR_3/XOR_0/NAND_2/w_32_0# comparator_0/XNOR_3/XOR_0/NAND_3/in2 0.03fF
C489 comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_32_0# 0.03fF
C490 gnd enableblock_1/enable1_1/AND_0/not_0/in 0.04fF
C491 comparator_0/A3 AND_2/in2 0.06fF
C492 comparator_0/A1 vdd 0.20fF
C493 enableblock_1/enable1_1/AND_0/NAND_0/w_32_0# enableblock_1/enable1_1/AND_0/not_0/in 0.03fF
C494 andblock_0/A3 gnd 0.10fF
C495 AND_1/NAND_0/w_32_0# AND_1/not_0/in 0.03fF
C496 addersubtractor_0/fulladder_2/OR_0/in2 gnd 0.36fF
C497 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_0_0# addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 0.03fF
C498 B2 B3 0.19fF
C499 comparator_0/XNOR_3/XOR_0/NAND_0/w_32_0# comparator_0/B0 0.06fF
C500 enableblock_0/B_out2 S0 0.06fF
C501 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_0_0# 0.05fF
C502 twotofourdecoder_0/AND_2/NAND_0/w_32_0# twotofourdecoder_0/AND_2/not_0/in 0.03fF
C503 B1 enableblock_2/enable1_1/AND_1/NAND_0/w_32_0# 0.06fF
C504 comparator_0/A0 vdd 0.26fF
C505 enableblock_0/enable1_1/AND_3/NAND_0/w_0_0# enableblock_0/enable1_1/AND_3/not_0/in 0.03fF
C506 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_0_0# vdd 0.05fF
C507 addersubtractor_0/fulladder_1/XOR_1/NAND_2/a_6_n14# addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 0.12fF
C508 addersubtractor_0/XOR_0/out addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_32_0# 0.06fF
C509 andblock_0/AND_0/NAND_0/w_0_0# vdd 0.05fF
C510 enableblock_0/enable1_1/AND_3/NAND_0/w_32_0# vdd 0.05fF
C511 gnd enableblock_1/enable1_1/AND_3/not_0/in 0.04fF
C512 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_32_0# 0.05fF
C513 addersubtractor_0/fulladder_1/XOR_1/NAND_2/a_6_n14# gnd 0.59fF
C514 comparator_0/AND_0/NAND_0/w_0_0# vdd 0.05fF
C515 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_32_0# 0.05fF
C516 addersubtractor_0/fulladder_0/OR_0/in1 vdd 0.12fF
C517 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_32_0# 0.05fF
C518 addersubtractor_0/fulladder_1/XOR_0/NAND_2/a_6_n14# gnd 0.59fF
C519 comparator_0/fourinputAND_1/fourinputNAND_0/w_63_0# comparator_0/XNOR_1/out 0.06fF
C520 enableblock_0/B_out2 addersubtractor_0/XOR_2/NAND_0/w_0_0# 0.06fF
C521 enableblock_0/B_out3 gnd 1.68fF
C522 addersubtractor_0/fulladder_1/XOR_0/NAND_2/a_6_n14# addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 0.12fF
C523 enableblock_2/enable1_0/AND_1/NAND_0/w_0_0# enableblock_2/En 0.06fF
C524 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_32_0# addersubtractor_0/XOR_3/out 0.06fF
C525 enableblock_0/enable1_1/AND_3/not_0/in vdd 0.29fF
C526 vdd addersubtractor_0/XOR_1/NAND_2/w_0_0# 0.05fF
C527 vdd addersubtractor_0/XOR_0/NAND_0/w_0_0# 0.05fF
C528 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_32_0# addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 0.03fF
C529 addersubtractor_0/fulladder_2/OR_0/in2 addersubtractor_0/fulladder_2/OR_0/NOR_0/w_32_0# 0.06fF
C530 twotofourdecoder_0/not_1/out twotofourdecoder_0/not_1/w_0_0# 0.03fF
C531 enableblock_2/enable1_0/AND_3/NAND_0/a_6_n14# gnd 0.57fF
C532 enableblock_2/enable1_0/AND_2/not_0/w_0_0# vdd 0.05fF
C533 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_0_0# adder3 0.03fF
C534 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_0_0# 0.05fF
C535 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_0/a_6_n14# 0.12fF
C536 twotofourdecoder_0/AND_1/NAND_0/w_32_0# twotofourdecoder_0/AND_1/not_0/in 0.03fF
C537 addersubtractor_0/fulladder_2/OR_0/in1 gnd 0.30fF
C538 comparator_0/fourinputAND_1/not_0/in comparator_0/XNOR_1/out 0.03fF
C539 gnd enableblock_1/enable1_1/AND_0/NAND_0/a_6_n14# 0.57fF
C540 vdd AND_2/not_0/w_0_0# 0.05fF
C541 enableblock_0/A_out2 gnd 0.92fF
C542 vdd addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# 0.21fF
C543 vdd addersubtractor_0/XOR_2/out 0.32fF
C544 addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_32_0# addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 0.03fF
C545 B3 S1 0.06fF
C546 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_0_0# addersubtractor_0/fulladder_3/XOR_1/in2 0.03fF
C547 A0 A1 0.20fF
C548 enableblock_2/enable1_0/AND_3/NAND_0/w_0_0# vdd 0.05fF
C549 enableblock_0/enable1_0/AND_0/NAND_0/w_32_0# OR_0/out 0.06fF
C550 andblock_0/AND_2/not_0/in vdd 0.29fF
C551 comparator_0/NOR_0/w_32_0# AND_1/in2 0.03fF
C552 vdd enableblock_1/enable1_1/AND_0/NAND_0/w_0_0# 0.05fF
C553 XOR_0/NAND_3/w_32_0# Carry 0.03fF
C554 andblock_0/AND_0/NAND_0/a_6_n14# andblock_0/AND_0/not_0/in 0.12fF
C555 comparator_0/XNOR_2/not_0/w_0_0# comparator_0/XNOR_2/not_0/in 0.06fF
C556 B3 enableblock_2/enable1_0/AND_1/NAND_0/w_32_0# 0.06fF
C557 comparator_0/A1 enableblock_1/enable1_1/AND_0/not_0/in 0.02fF
C558 addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_2/w_0_0# 0.06fF
C559 XOR_0/NAND_1/w_0_0# XOR_0/in1 0.06fF
C560 comparator_0/AND_0/out vdd 0.76fF
C561 enableblock_0/enable1_1/AND_1/NAND_0/w_32_0# enableblock_0/enable1_1/AND_1/not_0/in 0.03fF
C562 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_32_0# 0.03fF
C563 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/fulladder_1/AND_0/NAND_0/w_0_0# 0.03fF
C564 comparator_0/AND_0/out AND_2/in2 0.73fF
C565 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_0_0# 0.06fF
C566 comparator_0/XNOR_1/XOR_0/NAND_3/in1 gnd 0.11fF
C567 comparator_0/XNOR_1/XOR_0/NAND_1/w_0_0# vdd 0.05fF
C568 B0 A1 0.75fF
C569 XOR_0/NAND_2/in1 XOR_0/NAND_1/w_32_0# 0.06fF
C570 comparator_0/XNOR_3/not_0/w_0_0# comparator_0/XNOR_3/not_0/in 0.06fF
C571 andblock_0/AND_2/NAND_0/w_32_0# vdd 0.05fF
C572 andblock_0/A3 andblock_0/AND_0/NAND_0/w_0_0# 0.06fF
C573 gnd addersubtractor_0/XOR_2/NAND_3/in1 0.11fF
C574 and0 andblock_0/AND_3/not_0/in 0.02fF
C575 comparator_0/XNOR_0/XOR_0/NAND_3/in1 gnd 0.11fF
C576 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_0_0# 0.06fF
C577 andblock_0/A0 gnd 0.53fF
C578 comparator_0/XNOR_2/XOR_0/NAND_3/in1 gnd 0.11fF
C579 OR_0/NOR_0/w_32_0# OR_0/NOT_0/in 0.03fF
C580 enableblock_0/enable1_1/AND_3/not_0/w_0_0# enableblock_0/B_out0 0.03fF
C581 gnd AND_0/not_0/in 0.04fF
C582 addersubtractor_0/fulladder_0/OR_0/NOT_0/in gnd 0.60fF
C583 enableblock_0/enable1_1/AND_0/NAND_0/a_6_n14# A2 0.07fF
C584 addersubtractor_0/fulladder_0/OR_0/NOR_0/w_0_0# addersubtractor_0/fulladder_0/OR_0/in1 0.06fF
C585 comparator_0/XNOR_3/XOR_0/NAND_3/in1 gnd 0.11fF
C586 A3 gnd 0.32fF
C587 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/fulladder_2/AND_0/NAND_0/w_32_0# 0.03fF
C588 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 0.25fF
C589 AND_1/NAND_0/a_6_n14# AND_2/in2 0.07fF
C590 enableblock_0/B_out2 vdd 0.20fF
C591 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_0/a_6_n14# 0.12fF
C592 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 vdd 0.25fF
C593 enableblock_1/enable1_1/AND_0/NAND_0/w_0_0# enableblock_1/enable1_1/AND_0/not_0/in 0.03fF
C594 addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_32_0# addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 0.03fF
C595 addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_1/OR_0/NOR_0/w_0_0# 0.03fF
C596 twotofourdecoder_0/not_0/out S0 0.02fF
C597 twotofourdecoder_0/AND_2/NAND_0/w_32_0# vdd 0.05fF
C598 addersubtractor_0/fulladder_3/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_3/AND_1/not_0/in 0.03fF
C599 addersubtractor_0/XOR_0/NAND_1/w_32_0# addersubtractor_0/XOR_0/NAND_3/in1 0.03fF
C600 gnd addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 0.11fF
C601 B3 enableblock_2/En 0.13fF
C602 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_0_0# 0.05fF
C603 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_0_0# addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 0.03fF
C604 A3 OR_0/out 0.07fF
C605 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_32_0# addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 0.03fF
C606 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 gnd 0.11fF
C607 twotofourdecoder_0/AND_2/not_0/in vdd 0.29fF
C608 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_0_0# 0.05fF
C609 addersubtractor_0/fulladder_1/OR_0/NOT_0/in addersubtractor_0/fulladder_1/OR_0/NOR_0/w_32_0# 0.03fF
C610 S0 addersubtractor_0/XOR_1/NAND_0/w_32_0# 0.06fF
C611 comparator_0/threeinputAND_0/not_0/in comparator_0/threeinputAND_0/not_0/w_0_0# 0.06fF
C612 enableblock_0/B_out3 addersubtractor_0/XOR_2/out 0.11fF
C613 vdd S0 0.51fF
C614 addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_0_0# addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 0.03fF
C615 enableblock_0/A_out2 addersubtractor_0/XOR_0/NAND_0/w_0_0# 0.06fF
C616 comparator_0/XNOR_1/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_1/XOR_0/NAND_3/in2 0.06fF
C617 addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_0_0# 0.06fF
C618 comparator_0/fourinputAND_1/not_0/in comparator_0/XNOR_2/out 0.01fF
C619 enableblock_2/enable1_0/AND_2/NAND_0/w_32_0# enableblock_2/enable1_0/AND_2/not_0/in 0.03fF
C620 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_0_0# addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 0.03fF
C621 gnd addersubtractor_0/XOR_1/NAND_1/a_6_n14# 0.57fF
C622 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_0_0# vdd 0.05fF
C623 XOR_0/NAND_2/w_32_0# XOR_0/NAND_3/in2 0.03fF
C624 XOR_0/NAND_3/in2 vdd 0.25fF
C625 enableblock_0/B_out0 addersubtractor_0/XOR_3/NAND_0/w_0_0# 0.06fF
C626 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_0/AND_1/not_0/in 0.03fF
C627 addersubtractor_0/XOR_3/out addersubtractor_0/XOR_3/NAND_3/w_32_0# 0.03fF
C628 comparator_0/XNOR_1/not_0/in comparator_0/XNOR_1/XOR_0/NAND_3/a_6_n14# 0.12fF
C629 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_1/w_32_0# 0.06fF
C630 enableblock_2/enable1_1/AND_2/NAND_0/a_6_n14# enableblock_2/enable1_1/AND_2/not_0/in 0.12fF
C631 comparator_0/XNOR_3/out vdd 0.36fF
C632 comparator_0/fourinputAND_1/not_0/in gnd 0.01fF
C633 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_32_0# vdd 0.05fF
C634 comparator_0/XNOR_0/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_0/XOR_0/NAND_3/in2 0.06fF
C635 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# comparator_0/fourinputOR_0/not_0/in 0.04fF
C636 enableblock_1/enable1_0/AND_2/NAND_0/a_6_n14# gnd 0.57fF
C637 enableblock_1/enable1_0/AND_1/not_0/w_0_0# vdd 0.05fF
C638 addersubtractor_0/XOR_3/NAND_2/w_0_0# addersubtractor_0/XOR_3/NAND_3/in2 0.03fF
C639 vdd addersubtractor_0/XOR_2/NAND_0/w_0_0# 0.05fF
C640 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_0_0# 0.06fF
C641 comparator_0/threeinputAND_0/not_0/in comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# 0.11fF
C642 comparator_0/B2 gnd 0.22fF
C643 enableblock_1/enable1_1/AND_1/NAND_0/a_6_n14# enableblock_1/enable1_1/AND_1/not_0/in 0.12fF
C644 comparator_0/XNOR_0/not_0/in comparator_0/XNOR_0/XOR_0/NAND_3/a_6_n14# 0.12fF
C645 enableblock_1/enable1_0/AND_2/NAND_0/w_0_0# vdd 0.05fF
C646 OR_0/out enableblock_0/enable1_0/AND_3/NAND_0/w_0_0# 0.06fF
C647 enableblock_0/enable1_0/AND_2/NAND_0/w_0_0# A1 0.06fF
C648 addersubtractor_0/XOR_1/out addersubtractor_0/XOR_1/NAND_3/a_6_n14# 0.12fF
C649 comparator_0/XNOR_2/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_2/XOR_0/NAND_3/in2 0.06fF
C650 comparator_0/XNOR_1/XOR_0/NAND_2/in1 vdd 0.25fF
C651 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_100_0# comparator_0/fiveinputAND_0/not_0/in 0.03fF
C652 AND_2/in1 comparator_0/fourinputAND_1/not_0/in 0.02fF
C653 comparator_0/fourinputAND_0/not_0/in comparator_0/XNOR_0/out 0.01fF
C654 comparator_0/fourinputOR_0/in4 comparator_0/fiveinputAND_0/not_0/in 0.16fF
C655 comparator_0/fourinputOR_0/not_0/in comparator_0/fourinputOR_0/in2 0.11fF
C656 comparator_0/not_1/out vdd 0.07fF
C657 comparator_0/fourinputAND_0/fourinputNAND_0/w_100_0# vdd 0.05fF
C658 comparator_0/XNOR_2/not_0/in comparator_0/XNOR_2/XOR_0/NAND_3/a_6_n14# 0.12fF
C659 addersubtractor_0/XOR_0/out addersubtractor_0/XOR_0/NAND_3/a_6_n14# 0.12fF
C660 andblock_0/AND_0/NAND_0/w_32_0# andblock_0/AND_0/not_0/in 0.03fF
C661 comparator_0/not_3/out gnd 0.35fF
C662 comparator_0/XNOR_3/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_3/XOR_0/NAND_3/in2 0.06fF
C663 enableblock_1/enable1_0/AND_2/not_0/w_0_0# comparator_0/A2 0.03fF
C664 enableblock_0/B_out2 enableblock_0/B_out3 0.78fF
C665 twotofourdecoder_0/AND_0/NAND_0/w_32_0# vdd 0.05fF
C666 enableblock_2/enable1_0/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C667 enableblock_2/enable1_1/AND_0/NAND_0/w_32_0# enableblock_2/enable1_1/AND_0/not_0/in 0.03fF
C668 addersubtractor_0/fulladder_1/OR_0/NOT_0/in addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# 0.04fF
C669 enableblock_0/enable1_1/AND_3/NAND_0/a_6_n14# gnd 0.57fF
C670 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_0_0# 0.05fF
C671 enableblock_0/enable1_1/AND_2/not_0/w_0_0# vdd 0.05fF
C672 enableblock_1/enable1_0/AND_2/NAND_0/a_6_n14# enableblock_1/enable1_0/AND_2/not_0/in 0.12fF
C673 comparator_0/XNOR_3/not_0/in comparator_0/XNOR_3/XOR_0/NAND_3/a_6_n14# 0.12fF
C674 comparator_0/XNOR_0/not_0/w_0_0# comparator_0/XNOR_0/not_0/in 0.06fF
C675 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# gnd 0.35fF
C676 twotofourdecoder_0/AND_2/NAND_0/w_0_0# twotofourdecoder_0/AND_2/not_0/in 0.03fF
C677 vdd enableblock_1/enable1_0/AND_0/NAND_0/w_0_0# 0.05fF
C678 andblock_0/AND_3/NAND_0/w_0_0# vdd 0.05fF
C679 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_0_0# vdd 0.05fF
C680 addersubtractor_0/fulladder_0/XOR_1/in2 gnd 0.63fF
C681 comparator_0/fourinputAND_0/not_0/w_0_0# comparator_0/fourinputAND_0/not_0/in 0.06fF
C682 B3 A0 0.19fF
C683 andblock_0/AND_3/NAND_0/a_6_n14# gnd 0.57fF
C684 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_2/w_0_0# 0.06fF
C685 comparator_0/XNOR_1/XOR_0/NAND_1/w_0_0# comparator_0/XNOR_1/XOR_0/NAND_3/in1 0.03fF
C686 andblock_0/AND_1/not_0/w_0_0# vdd 0.05fF
C687 comparator_0/fourinputAND_1/fourinputNAND_0/w_32_0# vdd 0.05fF
C688 twotofourdecoder_0/not_0/out vdd 0.13fF
C689 twotofourdecoder_0/AND_3/not_0/w_0_0# twotofourdecoder_0/AND_3/not_0/in 0.06fF
C690 twotofourdecoder_0/AND_0/NAND_0/a_6_n14# twotofourdecoder_0/AND_0/not_0/in 0.12fF
C691 twotofourdecoder_0/AND_0/NAND_0/w_0_0# S0 0.06fF
C692 enableblock_0/enable1_1/AND_3/NAND_0/w_0_0# vdd 0.05fF
C693 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_32_0# 0.03fF
C694 addersubtractor_0/fulladder_1/XOR_1/NAND_3/a_6_n14# gnd 0.57fF
C695 andblock_0/AND_1/NAND_0/w_0_0# vdd 0.05fF
C696 enableblock_0/B_out3 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_0_0# 0.06fF
C697 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_32_0# 0.05fF
C698 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_1/w_32_0# 0.06fF
C699 comparator_0/B2 comparator_0/A1 0.76fF
C700 enableblock_2/enable1_0/AND_1/not_0/in gnd 0.04fF
C701 addersubtractor_0/fulladder_1/XOR_0/NAND_3/a_6_n14# gnd 0.57fF
C702 AND_2/in1 comparator_0/fourinputAND_1/not_0/w_0_0# 0.03fF
C703 gnd addersubtractor_0/XOR_3/out 0.56fF
C704 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_32_0# 0.05fF
C705 andblock_0/B3 enableblock_2/enable1_0/AND_1/not_0/in 0.02fF
C706 enableblock_0/B_out3 S0 0.06fF
C707 vdd vdd 0.05fF
C708 vdd addersubtractor_0/XOR_1/NAND_0/w_32_0# 0.05fF
C709 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_32_0# addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 0.06fF
C710 addersubtractor_0/fulladder_2/OR_0/NOT_0/in addersubtractor_0/fulladder_2/OR_0/NOT_0/w_0_0# 0.06fF
C711 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 gnd 0.15fF
C712 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_0_0# enableblock_0/A_out3 0.06fF
C713 XOR_0/NAND_2/w_32_0# vdd 0.05fF
C714 XOR_0/NAND_2/a_6_n14# gnd 0.59fF
C715 addersubtractor_0/fulladder_0/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_0/AND_1/not_0/in 0.06fF
C716 comparator_0/fourinputAND_0/fourinputNAND_0/w_32_0# comparator_0/A1 0.06fF
C717 twotofourdecoder_0/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C718 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_2/AND_1/not_0/in 0.03fF
C719 B2 B1 0.19fF
C720 B3 B0 0.19fF
C721 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_32_0# comparator_0/A0 0.06fF
C722 enableblock_0/enable1_1/AND_0/not_0/in vdd 0.29fF
C723 A2 gnd 0.32fF
C724 vdd addersubtractor_0/fulladder_3/OR_0/NOT_0/w_0_0# 0.05fF
C725 vdd addersubtractor_0/fulladder_2/AND_1/NAND_0/w_32_0# 0.05fF
C726 addersubtractor_0/fulladder_2/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C727 addersubtractor_0/fulladder_1/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_0/C 0.07fF
C728 comparator_0/XNOR_1/XOR_0/NAND_2/a_6_n14# comparator_0/XNOR_1/XOR_0/NAND_3/in2 0.12fF
C729 comparator_0/fiveinputAND_0/not_0/w_0_0# comparator_0/fiveinputAND_0/not_0/in 0.06fF
C730 enableblock_0/A_out2 S0 0.06fF
C731 addersubtractor_0/fulladder_2/XOR_1/NAND_0/a_6_n14# gnd 0.57fF
C732 AND_2/in1 AND_2/NAND_0/w_0_0# 0.06fF
C733 XOR_0/NAND_0/w_0_0# vdd 0.05fF
C734 enableblock_0/A_out0 addersubtractor_0/XOR_1/NAND_1/w_0_0# 0.06fF
C735 adder2 addersubtractor_0/fulladder_2/XOR_1/NAND_3/a_6_n14# 0.12fF
C736 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 0.06fF
C737 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_32_0# vdd 0.05fF
C738 vdd AND_2/in2 0.66fF
C739 S0 addersubtractor_0/XOR_2/NAND_2/w_32_0# 0.06fF
C740 comparator_0/NOR_0/a_13_6# AND_1/in2 0.04fF
C741 comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# vdd 0.21fF
C742 addersubtractor_0/fulladder_2/OR_0/NOT_0/w_0_0# addersubtractor_0/fulladder_2/C 0.03fF
C743 vdd addersubtractor_0/fulladder_1/C 0.18fF
C744 enableblock_0/enable1_0/AND_3/NAND_0/w_32_0# vdd 0.05fF
C745 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_3/a_6_n14# 0.12fF
C746 comparator_0/XNOR_0/XOR_0/NAND_2/a_6_n14# comparator_0/XNOR_0/XOR_0/NAND_3/in2 0.12fF
C747 A2 OR_0/out 0.07fF
C748 comparator_0/fourinputOR_0/fourinputNOR_0/w_97_0# vdd 0.03fF
C749 enableblock_0/enable1_0/AND_3/not_0/in vdd 0.29fF
C750 comparator_0/A0 enableblock_1/enable1_1/AND_2/not_0/w_0_0# 0.03fF
C751 vdd addersubtractor_0/XOR_2/NAND_3/in2 0.25fF
C752 greater comparator_0/fourinputOR_0/not_0/in 0.02fF
C753 enableblock_0/enable1_1/AND_0/not_0/w_0_0# vdd 0.05fF
C754 enableblock_0/enable1_1/AND_0/not_0/w_0_0# enableblock_0/enable1_1/AND_0/not_0/in 0.06fF
C755 enableblock_1/enable1_0/AND_0/NAND_0/a_6_n14# enableblock_1/enable1_0/AND_0/not_0/in 0.12fF
C756 comparator_0/XNOR_1/XOR_0/NAND_2/w_0_0# vdd 0.05fF
C757 comparator_0/fourinputOR_0/not_0/in comparator_0/fourinputOR_0/in3 0.15fF
C758 comparator_0/XNOR_2/XOR_0/NAND_2/a_6_n14# comparator_0/XNOR_2/XOR_0/NAND_3/in2 0.12fF
C759 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# comparator_0/A0 0.04fF
C760 B1 S1 0.06fF
C761 enableblock_2/enable1_1/AND_2/NAND_0/w_32_0# enableblock_2/En 0.06fF
C762 enableblock_0/enable1_0/AND_3/NAND_0/w_32_0# enableblock_0/enable1_0/AND_3/not_0/in 0.03fF
C763 comparator_0/XNOR_0/XOR_0/NAND_2/w_0_0# vdd 0.05fF
C764 addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/AND_0/not_0/in 0.02fF
C765 enableblock_2/enable1_1/AND_1/not_0/in vdd 0.29fF
C766 comparator_0/XNOR_2/XOR_0/NAND_2/w_0_0# vdd 0.05fF
C767 twotofourdecoder_0/AND_2/not_0/w_0_0# OR_0/in2 0.03fF
C768 vdd addersubtractor_0/XOR_3/NAND_1/w_0_0# 0.05fF
C769 addersubtractor_0/fulladder_1/AND_0/not_0/in gnd 0.04fF
C770 comparator_0/XNOR_3/XOR_0/NAND_2/a_6_n14# comparator_0/XNOR_3/XOR_0/NAND_3/in2 0.12fF
C771 twotofourdecoder_0/not_0/out twotofourdecoder_0/AND_2/NAND_0/w_0_0# 0.06fF
C772 vdd enableblock_1/enable1_1/AND_0/not_0/in 0.29fF
C773 enableblock_0/enable1_1/AND_3/NAND_0/a_6_n14# enableblock_0/enable1_1/AND_3/not_0/in 0.12fF
C774 addersubtractor_0/fulladder_2/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_2/AND_0/not_0/in 0.06fF
C775 addersubtractor_0/fulladder_1/XOR_0/NAND_0/a_6_n14# gnd 0.57fF
C776 twotofourdecoder_0/AND_2/NAND_0/a_6_n14# gnd 0.57fF
C777 andblock_0/A3 vdd 0.26fF
C778 vdd addersubtractor_0/fulladder_2/OR_0/in2 0.07fF
C779 vdd addersubtractor_0/fulladder_1/AND_1/not_0/w_0_0# 0.05fF
C780 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_1/AND_1/not_0/in 0.03fF
C781 XOR_0/NAND_0/w_32_0# OR_0/in1 0.06fF
C782 comparator_0/XNOR_3/XOR_0/NAND_2/w_0_0# vdd 0.05fF
C783 twotofourdecoder_0/AND_1/not_0/w_0_0# vdd 0.05fF
C784 gnd addersubtractor_0/XOR_0/NAND_0/a_6_n14# 0.57fF
C785 A3 S0 0.20fF
C786 vdd addersubtractor_0/XOR_2/NAND_1/w_32_0# 0.05fF
C787 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_0_0# 0.06fF
C788 addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_0_0# addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 0.03fF
C789 vdd enableblock_1/enable1_1/AND_3/NAND_0/w_32_0# 0.05fF
C790 twotofourdecoder_0/AND_1/not_0/w_0_0# AND_2/in2 0.03fF
C791 A0 enableblock_0/enable1_0/AND_0/NAND_0/a_6_n14# 0.07fF
C792 addersubtractor_0/fulladder_0/OR_0/NOR_0/w_0_0# vdd 0.05fF
C793 addersubtractor_0/fulladder_0/OR_0/NOT_0/w_0_0# addersubtractor_0/fulladder_0/C 0.03fF
C794 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_0_0# 0.05fF
C795 addersubtractor_0/fulladder_2/AND_1/not_0/in gnd 0.04fF
C796 twotofourdecoder_0/AND_2/NAND_0/w_0_0# vdd 0.05fF
C797 vdd addersubtractor_0/XOR_0/NAND_1/w_0_0# 0.05fF
C798 addersubtractor_0/fulladder_0/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_0/OR_0/in1 0.03fF
C799 andblock_0/AND_0/not_0/w_0_0# andblock_0/AND_0/not_0/in 0.06fF
C800 twotofourdecoder_0/AND_0/NAND_0/w_0_0# vdd 0.05fF
C801 vdd enableblock_1/enable1_1/AND_3/not_0/in 0.29fF
C802 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_0_0# addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 0.03fF
C803 enableblock_2/enable1_1/AND_0/not_0/in enableblock_2/enable1_1/AND_0/NAND_0/w_0_0# 0.03fF
C804 gnd addersubtractor_0/fulladder_3/OR_0/in2 0.36fF
C805 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_0_0# 0.05fF
C806 andblock_0/A2 gnd 0.36fF
C807 enableblock_0/enable1_0/AND_1/NAND_0/a_6_n14# enableblock_0/enable1_0/AND_1/not_0/in 0.12fF
C808 andblock_0/B3 andblock_0/A2 0.77fF
C809 gnd equal 0.08fF
C810 AND_0/in1 addersubtractor_0/fulladder_3/OR_0/NOT_0/in 0.02fF
C811 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_0_0# 0.05fF
C812 vdd enableblock_0/B_out3 0.30fF
C813 enableblock_0/enable1_0/AND_0/NAND_0/w_32_0# vdd 0.05fF
C814 enableblock_0/enable1_1/AND_0/not_0/in enableblock_0/B_out3 0.02fF
C815 addersubtractor_0/XOR_2/NAND_1/a_6_n14# addersubtractor_0/XOR_2/NAND_3/in1 0.12fF
C816 addersubtractor_0/fulladder_2/XOR_1/NAND_2/a_6_n14# addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 0.12fF
C817 comparator_0/fourinputOR_0/not_0/w_0_0# greater 0.03fF
C818 OR_0/in2 OR_0/NOR_0/w_32_0# 0.06fF
C819 enableblock_2/enable1_0/AND_2/NAND_0/w_0_0# enableblock_2/enable1_0/AND_2/not_0/in 0.03fF
C820 enableblock_0/A_out2 vdd 0.29fF
C821 A1 gnd 0.33fF
C822 vdd addersubtractor_0/fulladder_2/OR_0/in1 0.12fF
C823 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_0_0# S0 0.06fF
C824 XOR_0/NAND_3/w_32_0# XOR_0/NAND_3/in2 0.06fF
C825 addersubtractor_0/fulladder_2/XOR_0/NAND_2/a_6_n14# addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 0.12fF
C826 enableblock_2/enable1_0/AND_0/NAND_0/w_32_0# enableblock_2/enable1_0/AND_0/not_0/in 0.03fF
C827 comparator_0/AND_0/not_0/in gnd 0.04fF
C828 enableblock_2/enable1_0/AND_3/not_0/w_0_0# enableblock_2/enable1_0/AND_3/not_0/in 0.06fF
C829 AND_2/NAND_0/w_32_0# AND_2/not_0/in 0.03fF
C830 addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/AND_0/not_0/in 0.02fF
C831 andblock_0/AND_0/not_0/in gnd 0.04fF
C832 vdd addersubtractor_0/XOR_2/NAND_2/w_32_0# 0.05fF
C833 gnd addersubtractor_0/XOR_2/NAND_2/a_6_n14# 0.59fF
C834 Carry XOR_0/NAND_3/a_6_n14# 0.12fF
C835 enableblock_2/enable1_0/AND_0/not_0/in gnd 0.04fF
C836 B1 enableblock_2/En 0.13fF
C837 comparator_0/XNOR_1/not_0/in comparator_0/XNOR_1/out 0.02fF
C838 addersubtractor_0/XOR_2/out addersubtractor_0/XOR_2/NAND_3/w_32_0# 0.03fF
C839 addersubtractor_0/XOR_1/NAND_2/w_32_0# addersubtractor_0/XOR_1/NAND_3/in2 0.03fF
C840 OR_0/out A1 0.06fF
C841 andblock_0/A0 andblock_0/AND_3/NAND_0/w_0_0# 0.06fF
C842 enableblock_0/enable1_1/AND_0/not_0/w_0_0# enableblock_0/B_out3 0.03fF
C843 addersubtractor_0/XOR_3/NAND_2/in1 addersubtractor_0/XOR_3/NAND_2/w_0_0# 0.06fF
C844 enableblock_1/enable1_0/AND_3/not_0/in gnd 0.04fF
C845 gnd AND_0/NAND_0/a_6_n14# 0.57fF
C846 comparator_0/threeinputAND_0/not_0/w_0_0# comparator_0/fourinputOR_0/in2 0.03fF
C847 vdd addersubtractor_0/XOR_1/NAND_3/w_0_0# 0.05fF
C848 comparator_0/XNOR_1/XOR_0/NAND_3/in1 vdd 0.25fF
C849 A3 enableblock_1/enable1_0/AND_0/NAND_0/w_0_0# 0.06fF
C850 addersubtractor_0/fulladder_3/XOR_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 0.12fF
C851 addersubtractor_0/fulladder_1/AND_0/NAND_0/w_0_0# addersubtractor_0/XOR_1/out 0.06fF
C852 comparator_0/not_0/out comparator_0/not_0/w_0_0# 0.03fF
C853 comparator_0/B1 enableblock_1/enable1_1/AND_1/not_0/in 0.02fF
C854 addersubtractor_0/XOR_2/NAND_2/w_32_0# addersubtractor_0/XOR_2/NAND_3/in2 0.03fF
C855 vdd addersubtractor_0/XOR_2/NAND_3/in1 0.29fF
C856 addersubtractor_0/fulladder_1/AND_0/NAND_0/w_32_0# enableblock_0/A_out1 0.06fF
C857 comparator_0/XNOR_0/XOR_0/NAND_3/in1 vdd 0.25fF
C858 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/fulladder_2/AND_0/NAND_0/w_0_0# 0.03fF
C859 andblock_0/A0 vdd 0.20fF
C860 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_0_0# 0.06fF
C861 enableblock_1/enable1_1/AND_3/NAND_0/w_32_0# enableblock_1/enable1_1/AND_3/not_0/in 0.03fF
C862 enableblock_0/enable1_1/AND_1/not_0/in gnd 0.04fF
C863 addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_0/a_6_n14# 0.12fF
C864 comparator_0/XNOR_2/XOR_0/NAND_3/in1 vdd 0.25fF
C865 vdd AND_0/not_0/in 0.29fF
C866 andblock_0/AND_1/not_0/in and2 0.02fF
C867 addersubtractor_0/fulladder_0/OR_0/NOT_0/in vdd 0.11fF
C868 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_0_0# 0.06fF
C869 enableblock_1/enable1_1/AND_0/NAND_0/a_6_n14# enableblock_1/enable1_1/AND_0/not_0/in 0.12fF
C870 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_32_0# addersubtractor_0/XOR_2/out 0.06fF
C871 addersubtractor_0/fulladder_1/AND_1/not_0/in addersubtractor_0/fulladder_1/OR_0/in1 0.02fF
C872 comparator_0/XNOR_3/XOR_0/NAND_3/in1 vdd 0.25fF
C873 comparator_0/XNOR_1/not_0/w_0_0# comparator_0/XNOR_1/out 0.03fF
C874 addersubtractor_0/fulladder_0/XOR_1/in2 S0 0.06fF
C875 comparator_0/not_1/out comparator_0/B2 0.02fF
C876 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 0.15fF
C877 addersubtractor_0/fulladder_2/OR_0/NOT_0/in gnd 0.60fF
C878 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_0_0# 0.05fF
C879 comparator_0/fourinputOR_0/fourinputNOR_0/w_64_0# vdd 0.03fF
C880 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_1/a_6_n14# 0.12fF
C881 addersubtractor_0/fulladder_1/OR_0/NOR_0/w_0_0# addersubtractor_0/fulladder_1/OR_0/in1 0.06fF
C882 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_0_0# 0.03fF
C883 andblock_0/AND_0/not_0/w_0_0# and3 0.03fF
C884 addersubtractor_0/XOR_2/NAND_0/w_32_0# addersubtractor_0/XOR_2/NAND_2/in1 0.03fF
C885 enableblock_0/A_out2 addersubtractor_0/XOR_0/NAND_1/w_0_0# 0.06fF
C886 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 0.25fF
C887 enableblock_2/enable1_0/AND_2/not_0/w_0_0# andblock_0/A2 0.03fF
C888 comparator_0/fourinputAND_0/fourinputNAND_0/w_0_0# comparator_0/not_2/out 0.06fF
C889 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_1/a_6_n14# 0.12fF
C890 twotofourdecoder_0/not_1/w_0_0# vdd 0.05fF
C891 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 0.25fF
C892 addersubtractor_0/fulladder_0/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C893 addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_2/OR_0/NOR_0/w_0_0# 0.03fF
C894 addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/OR_0/NOR_0/w_32_0# 0.06fF
C895 addersubtractor_0/fulladder_0/AND_0/not_0/w_0_0# vdd 0.05fF
C896 XOR_0/NAND_3/a_6_n14# gnd 0.57fF
C897 XOR_0/NAND_3/w_32_0# vdd 0.05fF
C898 andblock_0/AND_0/NAND_0/w_0_0# andblock_0/AND_0/not_0/in 0.03fF
C899 comparator_0/fourinputAND_1/fourinputNAND_0/w_32_0# comparator_0/fourinputAND_1/not_0/in 0.03fF
C900 AND_2/not_0/w_0_0# equal 0.03fF
C901 addersubtractor_0/fulladder_0/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_0/AND_1/not_0/in 0.12fF
C902 A2 S0 0.18fF
C903 comparator_0/AND_0/NAND_0/w_0_0# comparator_0/AND_0/not_0/in 0.03fF
C904 gnd addersubtractor_0/fulladder_2/C 1.20fF
C905 addersubtractor_0/fulladder_0/AND_0/NAND_0/w_32_0# addersubtractor_0/fulladder_0/AND_0/not_0/in 0.03fF
C906 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_0_0# comparator_0/fiveinputAND_0/not_0/in 0.03fF
C907 comparator_0/fourinputAND_0/fourinputNAND_0/w_63_0# comparator_0/fourinputAND_0/not_0/in 0.03fF
C908 enableblock_0/enable1_0/AND_3/NAND_0/a_6_n14# gnd 0.57fF
C909 enableblock_0/enable1_0/AND_2/not_0/w_0_0# vdd 0.05fF
C910 comparator_0/XNOR_0/out comparator_0/A2 0.06fF
C911 comparator_0/fourinputAND_1/fourinputNAND_0/w_63_0# vdd 0.05fF
C912 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_0_0# vdd 0.05fF
C913 XOR_0/NAND_2/a_6_n14# XOR_0/NAND_3/in2 0.12fF
C914 comparator_0/not_1/w_0_0# comparator_0/not_1/out 0.03fF
C915 addersubtractor_0/fulladder_2/OR_0/NOT_0/in addersubtractor_0/fulladder_2/OR_0/NOR_0/w_32_0# 0.03fF
C916 enableblock_0/enable1_0/AND_1/not_0/w_0_0# enableblock_0/enable1_0/AND_1/not_0/in 0.06fF
C917 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_0_0# 0.03fF
C918 A0 B1 3.14fF
C919 addersubtractor_0/XOR_3/out addersubtractor_0/XOR_3/NAND_3/a_6_n14# 0.12fF
C920 vdd addersubtractor_0/fulladder_3/OR_0/NOR_0/w_32_0# 0.03fF
C921 and3 gnd 0.08fF
C922 lesser AND_1/not_0/in 0.02fF
C923 addersubtractor_0/XOR_2/NAND_1/w_32_0# addersubtractor_0/XOR_2/NAND_3/in1 0.03fF
C924 enableblock_0/enable1_0/AND_3/NAND_0/w_0_0# vdd 0.05fF
C925 comparator_0/fourinputAND_1/not_0/in vdd 1.27fF
C926 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_0_0# addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 0.03fF
C927 andblock_0/AND_1/NAND_0/a_6_n14# andblock_0/AND_1/not_0/in 0.12fF
C928 enableblock_1/enable1_0/AND_0/not_0/w_0_0# enableblock_1/enable1_0/AND_0/not_0/in 0.06fF
C929 A1 enableblock_1/enable1_1/AND_0/NAND_0/w_0_0# 0.06fF
C930 gnd AND_1/in2 0.95fF
C931 comparator_0/XNOR_0/out comparator_0/threeinputAND_0/threeinputNAND_0/w_63_0# 0.06fF
C932 comparator_0/not_2/out comparator_0/B1 0.02fF
C933 comparator_0/B2 vdd 0.30fF
C934 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_1/w_32_0# 0.06fF
C935 andblock_0/B0 enableblock_2/enable1_1/AND_3/not_0/in 0.02fF
C936 addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_1/w_32_0# 0.06fF
C937 addersubtractor_0/fulladder_1/OR_0/in2 addersubtractor_0/fulladder_1/OR_0/NOT_0/in 0.26fF
C938 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_32_0# vdd 0.05fF
C939 enableblock_1/enable1_0/AND_1/not_0/in enableblock_1/enable1_0/AND_1/NAND_0/w_0_0# 0.03fF
C940 comparator_0/threeinputAND_0/threeinputNAND_0/w_32_0# vdd 0.05fF
C941 comparator_0/not_2/w_0_0# comparator_0/not_2/out 0.03fF
C942 gnd addersubtractor_0/fulladder_3/AND_1/NAND_0/a_6_n14# 0.57fF
C943 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_0_0# adder0 0.03fF
C944 B0 B1 0.19fF
C945 comparator_0/XNOR_1/XOR_0/NAND_3/w_0_0# vdd 0.05fF
C946 comparator_0/XNOR_1/XOR_0/NAND_0/w_0_0# comparator_0/XNOR_1/XOR_0/NAND_2/in1 0.03fF
C947 comparator_0/XNOR_1/not_0/in gnd 0.03fF
C948 comparator_0/fourinputAND_0/fourinputNAND_0/w_32_0# vdd 0.05fF
C949 enableblock_1/enable1_0/AND_2/NAND_0/w_0_0# A2 0.06fF
C950 vdd AND_1/NAND_0/w_0_0# 0.05fF
C951 vdd addersubtractor_0/XOR_0/NAND_3/in2 0.25fF
C952 enableblock_0/enable1_1/AND_2/NAND_0/w_32_0# enableblock_0/enable1_1/AND_2/not_0/in 0.03fF
C953 addersubtractor_0/XOR_3/NAND_3/in1 addersubtractor_0/XOR_3/NAND_3/w_0_0# 0.06fF
C954 comparator_0/XNOR_2/out comparator_0/XNOR_2/not_0/in 0.02fF
C955 comparator_0/AND_0/out comparator_0/AND_0/not_0/in 0.02fF
C956 enableblock_2/enable1_1/AND_1/NAND_0/w_0_0# vdd 0.05fF
C957 enableblock_0/enable1_0/AND_0/not_0/in enableblock_0/A_out3 0.02fF
C958 comparator_0/fourinputOR_0/in4 gnd 0.21fF
C959 addersubtractor_0/XOR_3/NAND_0/w_0_0# addersubtractor_0/XOR_3/NAND_2/in1 0.03fF
C960 AND_2/in1 AND_1/in2 0.13fF
C961 comparator_0/XNOR_0/XOR_0/NAND_3/w_0_0# vdd 0.05fF
C962 comparator_0/XNOR_0/not_0/in gnd 0.03fF
C963 enableblock_0/enable1_0/AND_3/NAND_0/w_0_0# enableblock_0/enable1_0/AND_3/not_0/in 0.03fF
C964 AND_1/NAND_0/w_0_0# AND_2/in2 0.06fF
C965 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_0_0# addersubtractor_0/fulladder_0/XOR_1/in2 0.03fF
C966 comparator_0/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C967 enableblock_2/enable1_1/AND_3/not_0/w_0_0# vdd 0.05fF
C968 comparator_0/XNOR_0/out comparator_0/B1 0.06fF
C969 comparator_0/XNOR_2/not_0/in gnd 0.03fF
C970 XOR_0/NAND_2/in1 gnd 0.15fF
C971 comparator_0/XNOR_2/XOR_0/NAND_3/w_0_0# vdd 0.05fF
C972 comparator_0/not_3/out vdd 0.07fF
C973 twotofourdecoder_0/AND_2/NAND_0/a_6_n14# twotofourdecoder_0/AND_2/not_0/in 0.12fF
C974 gnd enableblock_1/enable1_1/AND_3/NAND_0/a_6_n14# 0.57fF
C975 vdd enableblock_1/enable1_1/AND_2/not_0/w_0_0# 0.05fF
C976 comparator_0/XNOR_0/out comparator_0/B0 0.06fF
C977 comparator_0/not_1/w_0_0# vdd 0.05fF
C978 comparator_0/XNOR_3/XOR_0/NAND_3/w_0_0# vdd 0.05fF
C979 comparator_0/XNOR_3/not_0/in gnd 0.03fF
C980 comparator_0/fourinputAND_1/not_0/w_0_0# vdd 0.05fF
C981 OR_0/NOR_0/a_13_6# vdd 0.21fF
C982 B3 gnd 0.91fF
C983 vdd adder0 0.25fF
C984 comparator_0/fourinputOR_0/in4 AND_2/in1 1.13fF
C985 vdd enableblock_1/enable1_1/AND_3/NAND_0/w_0_0# 0.05fF
C986 enableblock_0/enable1_0/AND_0/not_0/w_0_0# enableblock_0/A_out3 0.03fF
C987 addersubtractor_0/fulladder_0/XOR_1/in2 vdd 0.47fF
C988 andblock_0/AND_2/not_0/in andblock_0/AND_2/not_0/w_0_0# 0.06fF
C989 twotofourdecoder_0/AND_3/not_0/in gnd 0.04fF
C990 gnd enableblock_0/B_out1 1.65fF
C991 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_1/XOR_1/in2 0.06fF
C992 OR_0/in2 OR_0/in1 0.06fF
C993 comparator_0/XNOR_0/out comparator_0/XNOR_0/not_0/w_0_0# 0.03fF
C994 vdd addersubtractor_0/XOR_1/NAND_0/w_0_0# 0.05fF
C995 addersubtractor_0/fulladder_3/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_3/OR_0/in1 0.03fF
C996 enableblock_2/En enableblock_2/enable1_0/AND_2/NAND_0/w_32_0# 0.06fF
C997 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_0_0# enableblock_0/B_out1 0.06fF
C998 comparator_0/not_0/out comparator_0/B3 0.02fF
C999 enableblock_1/enable1_1/AND_3/NAND_0/w_0_0# AND_2/in2 0.06fF
C1000 vdd AND_2/NAND_0/w_0_0# 0.05fF
C1001 gnd addersubtractor_0/XOR_2/NAND_2/in1 0.15fF
C1002 addersubtractor_0/fulladder_2/OR_0/NOT_0/in addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# 0.04fF
C1003 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_0/XOR_1/in2 0.06fF
C1004 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_0_0# 0.05fF
C1005 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 gnd 0.15fF
C1006 addersubtractor_0/fulladder_0/AND_0/NAND_0/w_32_0# enableblock_0/A_out3 0.06fF
C1007 vdd addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# 0.21fF
C1008 gnd addersubtractor_0/fulladder_3/OR_0/in1 0.30fF
C1009 B3 OR_0/out 0.10fF
C1010 XOR_0/NAND_3/in1 XOR_0/NAND_1/w_0_0# 0.03fF
C1011 enableblock_2/enable1_0/AND_1/not_0/in vdd 0.29fF
C1012 vdd addersubtractor_0/XOR_3/out 0.32fF
C1013 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_0_0# 0.05fF
C1014 addersubtractor_0/fulladder_2/XOR_1/in2 gnd 0.63fF
C1015 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_0/C 0.06fF
C1016 addersubtractor_0/fulladder_1/AND_0/not_0/w_0_0# vdd 0.05fF
C1017 addersubtractor_0/fulladder_0/AND_1/not_0/w_0_0# vdd 0.05fF
C1018 enableblock_2/enable1_1/AND_1/NAND_0/w_0_0# enableblock_2/enable1_1/AND_1/not_0/in 0.03fF
C1019 enableblock_0/enable1_0/AND_2/not_0/in enableblock_0/A_out1 0.02fF
C1020 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 0.25fF
C1021 addersubtractor_0/fulladder_0/AND_0/NAND_0/a_6_n14# addersubtractor_0/XOR_0/out 0.07fF
C1022 comparator_0/XNOR_1/XOR_0/NAND_0/w_0_0# vdd 0.05fF
C1023 comparator_0/fourinputOR_0/not_0/in gnd 0.94fF
C1024 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_0_0# addersubtractor_0/fulladder_2/C 0.06fF
C1025 A1 S0 0.16fF
C1026 OR_0/out OR_0/NOT_0/w_0_0# 0.03fF
C1027 enableblock_2/enable1_1/AND_2/not_0/w_0_0# enableblock_2/enable1_1/AND_2/not_0/in 0.06fF
C1028 A2 AND_2/in2 0.06fF
C1029 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_32_0# addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 0.03fF
C1030 comparator_0/B3 comparator_0/XNOR_0/XOR_0/NAND_2/w_32_0# 0.06fF
C1031 vdd addersubtractor_0/XOR_2/NAND_3/w_32_0# 0.05fF
C1032 gnd addersubtractor_0/XOR_2/NAND_3/a_6_n14# 0.57fF
C1033 enableblock_1/enable1_1/AND_1/not_0/w_0_0# enableblock_1/enable1_1/AND_1/not_0/in 0.06fF
C1034 addersubtractor_0/fulladder_2/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_1/C 0.07fF
C1035 comparator_0/fourinputAND_0/not_0/w_0_0# comparator_0/fourinputOR_0/in3 0.03fF
C1036 addersubtractor_0/XOR_0/NAND_3/in1 addersubtractor_0/XOR_0/NAND_3/w_0_0# 0.06fF
C1037 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_0_0# addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 0.03fF
C1038 enableblock_0/B_out2 enableblock_0/enable1_1/AND_1/not_0/in 0.02fF
C1039 addersubtractor_0/fulladder_3/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_3/AND_1/not_0/in 0.03fF
C1040 vdd AND_1/NAND_0/w_32_0# 0.05fF
C1041 comparator_0/B1 comparator_0/XNOR_2/XOR_0/NAND_2/w_32_0# 0.06fF
C1042 enableblock_0/enable1_0/AND_3/not_0/w_0_0# enableblock_0/A_out0 0.03fF
C1043 A0 enableblock_2/enable1_1/AND_2/NAND_0/w_0_0# 0.06fF
C1044 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_0_0# addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 0.03fF
C1045 comparator_0/XNOR_0/XOR_0/NAND_0/w_32_0# vdd 0.05fF
C1046 addersubtractor_0/XOR_2/NAND_3/w_32_0# addersubtractor_0/XOR_2/NAND_3/in2 0.06fF
C1047 vdd enableblock_1/enable1_0/AND_1/NAND_0/w_32_0# 0.05fF
C1048 comparator_0/XNOR_2/XOR_0/NAND_0/w_32_0# vdd 0.05fF
C1049 enableblock_0/enable1_0/AND_1/NAND_0/w_32_0# enableblock_0/enable1_0/AND_1/not_0/in 0.03fF
C1050 comparator_0/B0 comparator_0/XNOR_3/XOR_0/NAND_2/w_32_0# 0.06fF
C1051 enableblock_0/enable1_1/AND_3/NAND_0/w_32_0# B3 0.06fF
C1052 comparator_0/B0 enableblock_1/enable1_1/AND_3/not_0/w_0_0# 0.03fF
C1053 enableblock_1/enable1_0/AND_2/not_0/w_0_0# enableblock_1/enable1_0/AND_2/not_0/in 0.06fF
C1054 enableblock_1/enable1_1/AND_3/NAND_0/w_0_0# enableblock_1/enable1_1/AND_3/not_0/in 0.03fF
C1055 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_0_0# 0.06fF
C1056 comparator_0/XNOR_3/XOR_0/NAND_0/w_32_0# vdd 0.05fF
C1057 vdd addersubtractor_0/fulladder_1/AND_0/not_0/in 0.29fF
C1058 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_32_0# vdd 0.05fF
C1059 addersubtractor_0/XOR_1/out gnd 0.56fF
C1060 enableblock_0/enable1_1/AND_1/NAND_0/w_0_0# OR_0/out 0.06fF
C1061 addersubtractor_0/fulladder_1/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_1/AND_1/not_0/in 0.12fF
C1062 enableblock_2/enable1_1/AND_0/NAND_0/w_32_0# vdd 0.05fF
C1063 enableblock_0/enable1_0/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C1064 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 0.11fF
C1065 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_0_0# 0.05fF
C1066 andblock_0/A2 andblock_0/AND_1/NAND_0/w_0_0# 0.06fF
C1067 twotofourdecoder_0/AND_3/NAND_0/w_0_0# twotofourdecoder_0/not_1/out 0.06fF
C1068 enableblock_2/enable1_1/AND_0/not_0/in andblock_0/A1 0.02fF
C1069 vdd addersubtractor_0/fulladder_2/AND_0/NAND_0/w_32_0# 0.05fF
C1070 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_32_0# addersubtractor_0/XOR_1/out 0.06fF
C1071 addersubtractor_0/XOR_0/NAND_3/in1 gnd 0.11fF
C1072 twotofourdecoder_0/AND_3/not_0/w_0_0# OR_0/in1 0.03fF
C1073 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 0.11fF
C1074 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_0_0# 0.05fF
C1075 comparator_0/A3 comparator_0/XNOR_0/XOR_0/NAND_1/w_0_0# 0.06fF
C1076 comparator_0/XNOR_1/XOR_0/NAND_3/in1 comparator_0/XNOR_1/XOR_0/NAND_3/w_0_0# 0.06fF
C1077 OR_0/out enableblock_0/enable1_1/AND_0/NAND_0/w_32_0# 0.06fF
C1078 vdd addersubtractor_0/fulladder_1/OR_0/NOT_0/w_0_0# 0.05fF
C1079 vdd addersubtractor_0/fulladder_2/AND_1/not_0/in 0.29fF
C1080 enableblock_2/enable1_1/AND_1/not_0/w_0_0# andblock_0/B1 0.03fF
C1081 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_2/AND_1/not_0/in 0.03fF
C1082 vdd enableblock_1/enable1_0/AND_0/NAND_0/w_32_0# 0.05fF
C1083 vdd addersubtractor_0/fulladder_3/OR_0/in2 0.07fF
C1084 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_0_0# 0.06fF
C1085 andblock_0/A2 vdd 0.20fF
C1086 comparator_0/fourinputAND_1/fourinputNAND_0/a_76_n14# comparator_0/XNOR_1/out 0.23fF
C1087 enableblock_2/enable1_0/AND_2/NAND_0/a_6_n14# enableblock_2/enable1_0/AND_2/not_0/in 0.12fF
C1088 enableblock_0/enable1_0/AND_1/not_0/in gnd 0.04fF
C1089 vdd addersubtractor_0/fulladder_2/OR_0/NOR_0/w_0_0# 0.05fF
C1090 enableblock_1/enable1_0/AND_0/NAND_0/w_32_0# AND_2/in2 0.06fF
C1091 vdd equal 0.09fF
C1092 addersubtractor_0/fulladder_1/OR_0/NOT_0/w_0_0# addersubtractor_0/fulladder_1/C 0.03fF
C1093 addersubtractor_0/fulladder_0/AND_1/NAND_0/a_6_n14# S0 0.07fF
C1094 OR_0/in1 OR_0/NOR_0/w_0_0# 0.06fF
C1095 comparator_0/A1 comparator_0/XNOR_2/XOR_0/NAND_1/w_0_0# 0.06fF
C1096 comparator_0/XNOR_0/XOR_0/NAND_3/in1 comparator_0/XNOR_0/XOR_0/NAND_3/w_0_0# 0.06fF
C1097 addersubtractor_0/XOR_0/NAND_3/in1 addersubtractor_0/XOR_0/NAND_1/a_6_n14# 0.12fF
C1098 vdd AND_0/NAND_0/w_0_0# 0.05fF
C1099 XOR_0/NAND_0/a_6_n14# gnd 0.57fF
C1100 OR_0/in2 OR_0/NOT_0/in 0.26fF
C1101 enableblock_2/enable1_1/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C1102 enableblock_2/enable1_1/AND_0/not_0/w_0_0# andblock_0/A1 0.03fF
C1103 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/fulladder_1/AND_0/NAND_0/a_6_n14# 0.12fF
C1104 comparator_0/A0 comparator_0/XNOR_3/XOR_0/NAND_1/w_0_0# 0.06fF
C1105 comparator_0/XNOR_2/XOR_0/NAND_3/in1 comparator_0/XNOR_2/XOR_0/NAND_3/w_0_0# 0.06fF
C1106 comparator_0/AND_0/not_0/in vdd 0.29fF
C1107 A1 AND_2/in2 0.06fF
C1108 andblock_0/AND_0/not_0/in vdd 0.29fF
C1109 enableblock_2/enable1_0/AND_0/not_0/in vdd 0.29fF
C1110 enableblock_1/enable1_0/AND_3/NAND_0/w_32_0# vdd 0.05fF
C1111 addersubtractor_0/XOR_2/out addersubtractor_0/XOR_2/NAND_3/a_6_n14# 0.12fF
C1112 comparator_0/fourinputAND_1/fourinputNAND_0/w_63_0# comparator_0/fourinputAND_1/not_0/in 0.03fF
C1113 andblock_0/A0 andblock_0/AND_3/NAND_0/a_6_n14# 0.02fF
C1114 comparator_0/fourinputOR_0/not_0/in comparator_0/AND_0/out 0.67fF
C1115 enableblock_1/enable1_0/AND_3/not_0/in vdd 0.29fF
C1116 comparator_0/XNOR_3/XOR_0/NAND_3/in1 comparator_0/XNOR_3/XOR_0/NAND_3/w_0_0# 0.06fF
C1117 A3 enableblock_2/enable1_0/AND_0/NAND_0/a_6_n14# 0.07fF
C1118 comparator_0/XNOR_0/out comparator_0/XNOR_1/out 1.10fF
C1119 enableblock_2/enable1_1/AND_2/not_0/in gnd 0.04fF
C1120 enableblock_0/enable1_1/AND_2/NAND_0/w_0_0# enableblock_0/enable1_1/AND_2/not_0/in 0.03fF
C1121 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_32_0# 0.05fF
C1122 addersubtractor_0/fulladder_0/XOR_1/NAND_1/a_6_n14# gnd 0.57fF
C1123 gnd enableblock_1/enable1_1/AND_1/not_0/in 0.04fF
C1124 addersubtractor_0/XOR_3/NAND_1/w_32_0# addersubtractor_0/XOR_3/NAND_3/in1 0.03fF
C1125 addersubtractor_0/XOR_2/NAND_2/a_6_n14# addersubtractor_0/XOR_2/NAND_3/in2 0.12fF
C1126 enableblock_0/enable1_1/AND_3/not_0/w_0_0# enableblock_0/enable1_1/AND_3/not_0/in 0.06fF
C1127 addersubtractor_0/fulladder_0/XOR_0/NAND_1/a_6_n14# gnd 0.57fF
C1128 enableblock_2/enable1_0/AND_0/not_0/w_0_0# vdd 0.05fF
C1129 addersubtractor_0/XOR_1/out addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_32_0# 0.06fF
C1130 twotofourdecoder_0/AND_0/not_0/w_0_0# twotofourdecoder_0/AND_0/not_0/in 0.06fF
C1131 enableblock_0/enable1_1/AND_1/not_0/in vdd 0.29fF
C1132 addersubtractor_0/fulladder_3/AND_0/NAND_0/w_32_0# addersubtractor_0/fulladder_3/AND_0/not_0/in 0.03fF
C1133 andblock_0/AND_2/not_0/w_0_0# vdd 0.05fF
C1134 addersubtractor_0/XOR_3/NAND_2/in1 addersubtractor_0/XOR_3/NAND_0/a_6_n14# 0.12fF
C1135 addersubtractor_0/fulladder_2/AND_0/NAND_0/w_0_0# addersubtractor_0/XOR_2/out 0.06fF
C1136 addersubtractor_0/fulladder_2/AND_0/NAND_0/w_32_0# enableblock_0/B_out3 0.06fF
C1137 twotofourdecoder_0/AND_3/NAND_0/w_32_0# S0 0.06fF
C1138 comparator_0/not_3/w_0_0# comparator_0/B0 0.06fF
C1139 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_0/a_6_n14# 0.12fF
C1140 B3 S0 0.17fF
C1141 comparator_0/fourinputOR_0/in4 comparator_0/XNOR_3/out 0.06fF
C1142 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_0_0# 0.06fF
C1143 B2 S1 0.06fF
C1144 A2 A3 0.19fF
C1145 andblock_0/A1 gnd 0.22fF
C1146 S0 enableblock_0/B_out1 0.06fF
C1147 enableblock_2/enable1_0/AND_1/NAND_0/w_0_0# vdd 0.05fF
C1148 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 0.25fF
C1149 vdd addersubtractor_0/fulladder_2/OR_0/NOT_0/in 0.11fF
C1150 gnd lesser 0.08fF
C1151 addersubtractor_0/fulladder_0/OR_0/in2 gnd 0.36fF
C1152 comparator_0/threeinputAND_0/not_0/in comparator_0/fourinputOR_0/in2 0.02fF
C1153 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_32_0# 0.06fF
C1154 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_0_0# 0.06fF
C1155 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_32_0# 0.06fF
C1156 addersubtractor_0/fulladder_2/AND_1/not_0/in addersubtractor_0/fulladder_2/OR_0/in1 0.02fF
C1157 comparator_0/XNOR_3/out comparator_0/XNOR_3/not_0/in 0.02fF
C1158 comparator_0/fourinputAND_1/not_0/w_0_0# comparator_0/fourinputAND_1/not_0/in 0.06fF
C1159 twotofourdecoder_0/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C1160 enableblock_2/enable1_0/AND_3/not_0/w_0_0# vdd 0.05fF
C1161 andblock_0/A3 enableblock_2/enable1_0/AND_0/not_0/in 0.02fF
C1162 enableblock_2/enable1_1/AND_0/NAND_0/w_0_0# vdd 0.05fF
C1163 enableblock_1/enable1_0/AND_1/not_0/in comparator_0/B3 0.02fF
C1164 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_0/a_6_n14# 0.57fF
C1165 comparator_0/not_1/w_0_0# comparator_0/B2 0.06fF
C1166 lesser AND_1/not_0/w_0_0# 0.03fF
C1167 comparator_0/fourinputAND_0/fourinputNAND_0/w_0_0# comparator_0/fourinputAND_0/not_0/in 0.03fF
C1168 andblock_0/AND_3/not_0/in gnd 0.04fF
C1169 addersubtractor_0/fulladder_2/OR_0/NOR_0/w_0_0# addersubtractor_0/fulladder_2/OR_0/in1 0.06fF
C1170 comparator_0/threeinputAND_0/not_0/in comparator_0/threeinputAND_0/threeinputNAND_0/w_0_0# 0.03fF
C1171 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_0/a_6_n14# 0.12fF
C1172 vdd addersubtractor_0/fulladder_2/C 0.18fF
C1173 addersubtractor_0/fulladder_0/AND_0/NAND_0/a_6_n14# addersubtractor_0/fulladder_0/AND_0/not_0/in 0.12fF
C1174 addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_0/w_0_0# 0.03fF
C1175 addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_3/OR_0/NOR_0/w_32_0# 0.03fF
C1176 B1 gnd 0.86fF
C1177 comparator_0/fourinputAND_1/fourinputNAND_0/a_76_n14# gnd 0.04fF
C1178 enableblock_0/enable1_0/AND_0/NAND_0/w_0_0# enableblock_0/enable1_0/AND_0/not_0/in 0.03fF
C1179 andblock_0/AND_3/NAND_0/w_32_0# vdd 0.05fF
C1180 comparator_0/not_2/out comparator_0/XNOR_2/out 0.06fF
C1181 comparator_0/XNOR_1/XOR_0/NAND_0/a_6_n14# gnd 0.57fF
C1182 comparator_0/threeinputAND_0/not_0/in comparator_0/threeinputAND_0/threeinputNAND_0/w_63_0# 0.03fF
C1183 A1 enableblock_1/enable1_1/AND_0/NAND_0/a_6_n14# 0.07fF
C1184 addersubtractor_0/XOR_1/NAND_2/w_0_0# addersubtractor_0/XOR_1/NAND_3/in2 0.03fF
C1185 and3 vdd 0.20fF
C1186 comparator_0/fourinputAND_0/fourinputNAND_0/a_45_n14# comparator_0/fourinputAND_0/fourinputNAND_0/a_76_n14# 0.04fF
C1187 enableblock_2/enable1_0/AND_0/not_0/w_0_0# andblock_0/A3 0.03fF
C1188 comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# gnd 0.47fF
C1189 comparator_0/XNOR_1/XOR_0/NAND_3/in2 gnd 0.07fF
C1190 comparator_0/not_2/out gnd 0.08fF
C1191 OR_0/out B1 0.07fF
C1192 enableblock_0/enable1_0/AND_0/not_0/in gnd 0.04fF
C1193 vdd addersubtractor_0/XOR_0/NAND_3/w_32_0# 0.05fF
C1194 gnd addersubtractor_0/XOR_0/NAND_3/a_6_n14# 0.57fF
C1195 vdd AND_1/in2 0.37fF
C1196 comparator_0/not_3/out comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# 0.10fF
C1197 AND_1/in2 AND_2/in2 0.06fF
C1198 comparator_0/XNOR_0/XOR_0/NAND_3/in2 gnd 0.07fF
C1199 enableblock_0/enable1_0/AND_3/NAND_0/a_6_n14# enableblock_0/enable1_0/AND_3/not_0/in 0.12fF
C1200 addersubtractor_0/XOR_3/NAND_1/w_32_0# addersubtractor_0/XOR_3/NAND_2/in1 0.06fF
C1201 andblock_0/AND_2/not_0/in andblock_0/AND_2/NAND_0/w_0_0# 0.03fF
C1202 gnd addersubtractor_0/XOR_1/NAND_2/in1 0.15fF
C1203 comparator_0/XNOR_0/out comparator_0/XNOR_2/out 0.51fF
C1204 comparator_0/XNOR_1/not_0/in vdd 0.25fF
C1205 andblock_0/B0 gnd 0.28fF
C1206 addersubtractor_0/fulladder_3/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_3/XOR_1/in2 0.06fF
C1207 andblock_0/AND_3/not_0/w_0_0# vdd 0.05fF
C1208 XOR_0/in1 gnd 0.88fF
C1209 comparator_0/XNOR_2/XOR_0/NAND_3/in2 gnd 0.07fF
C1210 addersubtractor_0/fulladder_2/OR_0/in2 addersubtractor_0/fulladder_2/OR_0/NOT_0/in 0.26fF
C1211 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_100_0# vdd 0.05fF
C1212 enableblock_2/En twotofourdecoder_0/AND_0/not_0/in 0.11fF
C1213 enableblock_0/enable1_1/AND_2/not_0/w_0_0# enableblock_0/B_out1 0.03fF
C1214 comparator_0/XNOR_0/not_0/in vdd 0.25fF
C1215 comparator_0/fourinputOR_0/in4 vdd 0.93fF
C1216 B2 enableblock_2/En 0.13fF
C1217 addersubtractor_0/XOR_1/NAND_1/w_32_0# addersubtractor_0/XOR_1/NAND_3/in1 0.03fF
C1218 gnd addersubtractor_0/XOR_1/NAND_0/a_6_n14# 0.57fF
C1219 comparator_0/XNOR_3/XOR_0/NAND_3/in2 gnd 0.07fF
C1220 comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# comparator_0/threeinputAND_0/threeinputNAND_0/a_45_n14# 0.04fF
C1221 comparator_0/XNOR_0/out gnd 0.98fF
C1222 addersubtractor_0/fulladder_3/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_3/AND_1/not_0/in 0.06fF
C1223 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_0_0# adder1 0.03fF
C1224 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 0.25fF
C1225 comparator_0/XNOR_2/not_0/in vdd 0.25fF
C1226 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_113_n14# gnd 0.04fF
C1227 XOR_0/NAND_2/in1 vdd 0.25fF
C1228 AND_0/not_0/in AND_0/NAND_0/w_0_0# 0.03fF
C1229 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 vdd 0.25fF
C1230 comparator_0/fourinputOR_0/in3 comparator_0/fourinputAND_0/not_0/in 0.02fF
C1231 gnd addersubtractor_0/fulladder_3/AND_1/not_0/in 0.04fF
C1232 addersubtractor_0/XOR_3/NAND_0/w_32_0# addersubtractor_0/XOR_3/NAND_2/in1 0.03fF
C1233 vdd addersubtractor_0/fulladder_2/AND_0/not_0/w_0_0# 0.05fF
C1234 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_0_0# addersubtractor_0/fulladder_1/XOR_1/in2 0.03fF
C1235 addersubtractor_0/fulladder_0/XOR_0/NAND_0/a_6_n14# gnd 0.57fF
C1236 XOR_0/NAND_2/in1 XOR_0/NAND_0/w_0_0# 0.03fF
C1237 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_0/w_0_0# 0.03fF
C1238 twotofourdecoder_0/AND_3/NAND_0/w_32_0# vdd 0.05fF
C1239 vdd addersubtractor_0/XOR_1/NAND_1/w_0_0# 0.05fF
C1240 comparator_0/XNOR_3/not_0/in vdd 0.25fF
C1241 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# 0.04fF
C1242 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_0_0# 0.05fF
C1243 addersubtractor_0/fulladder_0/XOR_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 0.12fF
C1244 A3 A1 0.19fF
C1245 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_0_0# 0.05fF
C1246 addersubtractor_0/fulladder_0/C gnd 1.14fF
C1247 comparator_0/fourinputOR_0/in4 comparator_0/fourinputOR_0/fourinputNOR_0/w_97_0# 0.06fF
C1248 twotofourdecoder_0/AND_3/not_0/in vdd 0.29fF
C1249 enableblock_2/En twotofourdecoder_0/AND_0/not_0/w_0_0# 0.03fF
C1250 B3 AND_2/in2 0.06fF
C1251 vdd enableblock_0/B_out1 0.29fF
C1252 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_0_0# vdd 0.05fF
C1253 twotofourdecoder_0/AND_1/NAND_0/w_32_0# twotofourdecoder_0/not_0/out 0.06fF
C1254 vdd addersubtractor_0/XOR_2/NAND_2/in1 0.25fF
C1255 enableblock_0/A_out3 addersubtractor_0/XOR_0/out 0.11fF
C1256 OR_0/NOT_0/w_0_0# vdd 0.05fF
C1257 comparator_0/XNOR_1/not_0/w_0_0# vdd 0.05fF
C1258 vdd addersubtractor_0/XOR_3/NAND_2/w_0_0# 0.05fF
C1259 vdd adder2 0.25fF
C1260 vdd addersubtractor_0/fulladder_3/OR_0/in1 0.12fF
C1261 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 0.25fF
C1262 XOR_0/NAND_3/in1 XOR_0/NAND_1/w_32_0# 0.03fF
C1263 comparator_0/not_0/out gnd 0.08fF
C1264 vdd addersubtractor_0/fulladder_2/XOR_1/in2 0.47fF
C1265 vdd addersubtractor_0/fulladder_1/OR_0/NOR_0/w_32_0# 0.03fF
C1266 enableblock_2/En S1 0.07fF
C1267 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_2/XOR_1/in2 0.06fF
C1268 AND_0/NAND_0/a_6_n14# AND_0/not_0/in 0.12fF
C1269 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_32_0# 0.06fF
C1270 twotofourdecoder_0/AND_1/NAND_0/w_32_0# vdd 0.05fF
C1271 comparator_0/fourinputAND_0/fourinputNAND_0/a_45_n14# comparator_0/A1 0.21fF
C1272 enableblock_0/enable1_0/AND_1/NAND_0/w_0_0# OR_0/out 0.06fF
C1273 addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/OR_0/NOR_0/w_32_0# 0.06fF
C1274 enableblock_0/enable1_1/AND_1/NAND_0/w_32_0# B2 0.06fF
C1275 OR_0/out AND_0/NAND_0/w_32_0# 0.06fF
C1276 comparator_0/XNOR_0/out comparator_0/A3 0.01fF
C1277 comparator_0/fourinputOR_0/not_0/in vdd 0.10fF
C1278 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 gnd 0.15fF
C1279 comparator_0/fiveinputAND_0/not_0/w_0_0# vdd 0.05fF
C1280 enableblock_1/enable1_0/AND_3/NAND_0/a_6_n14# gnd 0.57fF
C1281 enableblock_1/enable1_0/AND_2/not_0/w_0_0# vdd 0.05fF
C1282 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_1/C 0.06fF
C1283 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_1/a_6_n14# 0.12fF
C1284 comparator_0/XNOR_0/out comparator_0/A1 0.06fF
C1285 gnd addersubtractor_0/XOR_3/NAND_0/a_6_n14# 0.57fF
C1286 enableblock_0/B_out2 addersubtractor_0/XOR_2/NAND_1/w_0_0# 0.06fF
C1287 enableblock_1/enable1_0/AND_3/NAND_0/w_0_0# vdd 0.05fF
C1288 comparator_0/XNOR_0/out comparator_0/A0 0.06fF
C1289 addersubtractor_0/fulladder_1/OR_0/in2 gnd 0.36fF
C1290 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_1/a_6_n14# 0.12fF
C1291 comparator_0/XNOR_0/XOR_0/NAND_1/w_0_0# vdd 0.05fF
C1292 XOR_0/NAND_3/in1 XOR_0/NAND_3/w_0_0# 0.06fF
C1293 addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_32_0# addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 0.03fF
C1294 addersubtractor_0/fulladder_2/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_2/OR_0/in2 0.03fF
C1295 enableblock_1/enable1_0/AND_3/NAND_0/w_0_0# AND_2/in2 0.06fF
C1296 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_0/w_0_0# 0.03fF
C1297 comparator_0/fourinputOR_0/not_0/in comparator_0/fourinputOR_0/fourinputNOR_0/w_97_0# 0.03fF
C1298 addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_2/w_0_0# 0.06fF
C1299 comparator_0/XNOR_2/XOR_0/NAND_1/w_0_0# vdd 0.05fF
C1300 twotofourdecoder_0/AND_1/NAND_0/w_0_0# twotofourdecoder_0/AND_1/not_0/in 0.03fF
C1301 B2 A0 0.19fF
C1302 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_0_0# addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 0.03fF
C1303 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_32_0# addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 0.03fF
C1304 enableblock_1/enable1_1/AND_3/NAND_0/a_6_n14# enableblock_1/enable1_1/AND_3/not_0/in 0.12fF
C1305 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_32_0# 0.05fF
C1306 addersubtractor_0/fulladder_0/XOR_1/NAND_2/a_6_n14# gnd 0.59fF
C1307 twotofourdecoder_0/AND_2/not_0/w_0_0# twotofourdecoder_0/AND_2/not_0/in 0.06fF
C1308 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_32_0# 0.05fF
C1309 comparator_0/XNOR_3/XOR_0/NAND_1/w_0_0# vdd 0.05fF
C1310 enableblock_0/enable1_1/AND_1/NAND_0/w_0_0# vdd 0.05fF
C1311 addersubtractor_0/XOR_1/NAND_2/a_6_n14# addersubtractor_0/XOR_1/NAND_3/in2 0.12fF
C1312 addersubtractor_0/fulladder_1/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_1/AND_0/not_0/in 0.06fF
C1313 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_32_0# vdd 0.05fF
C1314 addersubtractor_0/fulladder_0/XOR_0/NAND_2/a_6_n14# gnd 0.59fF
C1315 addersubtractor_0/XOR_2/NAND_1/w_32_0# addersubtractor_0/XOR_2/NAND_2/in1 0.06fF
C1316 addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_0_0# addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 0.03fF
C1317 enableblock_0/A_out1 gnd 1.72fF
C1318 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_1/w_32_0# 0.06fF
C1319 vdd addersubtractor_0/fulladder_2/AND_0/NAND_0/w_0_0# 0.05fF
C1320 enableblock_0/enable1_1/AND_3/not_0/w_0_0# vdd 0.05fF
C1321 twotofourdecoder_0/AND_3/NAND_0/a_6_n14# twotofourdecoder_0/not_1/out 0.07fF
C1322 vdd enableblock_0/enable1_1/AND_0/NAND_0/w_32_0# 0.05fF
C1323 gnd enableblock_1/enable1_0/AND_0/NAND_0/a_6_n14# 0.57fF
C1324 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_32_0# addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 0.03fF
C1325 enableblock_0/enable1_1/AND_0/not_0/in enableblock_0/enable1_1/AND_0/NAND_0/w_32_0# 0.03fF
C1326 enableblock_1/enable1_0/AND_3/not_0/in comparator_0/B2 0.02fF
C1327 gnd addersubtractor_0/fulladder_3/OR_0/NOT_0/in 0.60fF
C1328 addersubtractor_0/fulladder_1/OR_0/in1 gnd 0.30fF
C1329 vdd addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# 0.21fF
C1330 B2 B0 0.19fF
C1331 vdd addersubtractor_0/XOR_1/out 0.32fF
C1332 comparator_0/fourinputOR_0/not_0/w_0_0# vdd 0.05fF
C1333 S1 twotofourdecoder_0/AND_1/NAND_0/w_0_0# 0.06fF
C1334 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 0.25fF
C1335 OR_0/in1 gnd 0.11fF
C1336 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_0_0# 0.06fF
C1337 enableblock_2/enable1_0/AND_2/not_0/in gnd 0.04fF
C1338 vdd addersubtractor_0/XOR_0/NAND_3/in1 0.25fF
C1339 comparator_0/not_0/out comparator_0/AND_0/NAND_0/w_0_0# 0.06fF
C1340 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_32_0# adder3 0.03fF
C1341 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 0.25fF
C1342 comparator_0/AND_0/out comparator_0/XNOR_0/out 0.06fF
C1343 comparator_0/not_0/w_0_0# comparator_0/B3 0.06fF
C1344 gnd AND_2/not_0/in 0.04fF
C1345 addersubtractor_0/fulladder_2/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_2/AND_1/not_0/in 0.12fF
C1346 A0 S1 0.06fF
C1347 comparator_0/A1 enableblock_1/enable1_1/AND_0/not_0/w_0_0# 0.03fF
C1348 twotofourdecoder_0/AND_0/NAND_0/a_6_n14# S0 0.11fF
C1349 enableblock_2/enable1_0/AND_0/NAND_0/a_6_n14# enableblock_2/enable1_0/AND_0/not_0/in 0.12fF
C1350 and1 gnd 0.08fF
C1351 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_3/XOR_1/in2 0.03fF
C1352 OR_0/out OR_0/in1 0.06fF
C1353 enableblock_0/enable1_0/AND_1/not_0/in vdd 0.29fF
C1354 comparator_0/fourinputAND_0/fourinputNAND_0/w_63_0# comparator_0/XNOR_1/out 0.06fF
C1355 comparator_0/AND_0/NAND_0/w_32_0# comparator_0/A3 0.06fF
C1356 andblock_0/B2 enableblock_2/enable1_0/AND_3/not_0/in 0.02fF
C1357 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_32_0# addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 0.06fF
C1358 B1 S0 0.16fF
C1359 vdd addersubtractor_0/XOR_3/NAND_0/w_0_0# 0.05fF
C1360 A2 A1 0.19fF
C1361 B0 S1 0.06fF
C1362 comparator_0/fourinputAND_0/not_0/in comparator_0/XNOR_1/out 0.03fF
C1363 enableblock_0/enable1_0/AND_2/NAND_0/w_32_0# enableblock_0/enable1_0/AND_2/not_0/in 0.03fF
C1364 comparator_0/XNOR_1/XOR_0/NAND_1/w_32_0# vdd 0.05fF
C1365 comparator_0/XNOR_1/XOR_0/NAND_1/a_6_n14# gnd 0.57fF
C1366 addersubtractor_0/fulladder_1/AND_0/NAND_0/a_6_n14# addersubtractor_0/XOR_1/out 0.07fF
C1367 andblock_0/AND_2/NAND_0/w_0_0# vdd 0.05fF
C1368 vdd addersubtractor_0/XOR_1/NAND_3/in2 0.25fF
C1369 comparator_0/XNOR_0/XOR_0/NAND_1/a_6_n14# gnd 0.57fF
C1370 enableblock_2/enable1_0/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C1371 enableblock_0/enable1_1/AND_2/NAND_0/a_6_n14# enableblock_0/enable1_1/AND_2/not_0/in 0.12fF
C1372 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/fulladder_2/AND_0/NAND_0/a_6_n14# 0.12fF
C1373 enableblock_2/enable1_1/AND_2/NAND_0/w_32_0# vdd 0.05fF
C1374 comparator_0/XNOR_2/XOR_0/NAND_1/a_6_n14# gnd 0.57fF
C1375 vdd enableblock_1/enable1_1/AND_1/NAND_0/w_32_0# 0.05fF
C1376 A3 B3 0.23fF
C1377 enableblock_2/enable1_1/AND_2/not_0/in vdd 0.29fF
C1378 comparator_0/XNOR_3/XOR_0/NAND_1/a_6_n14# gnd 0.57fF
C1379 comparator_0/fourinputAND_1/fourinputNAND_0/a_45_n14# comparator_0/fourinputAND_1/fourinputNAND_0/a_76_n14# 0.04fF
C1380 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 gnd 0.11fF
C1381 and2 gnd 0.08fF
C1382 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_0_0# 0.05fF
C1383 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_32_0# 0.06fF
C1384 vdd enableblock_1/enable1_1/AND_1/not_0/in 0.29fF
C1385 addersubtractor_0/XOR_3/NAND_1/a_6_n14# addersubtractor_0/XOR_3/NAND_3/in1 0.12fF
C1386 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_1/w_32_0# 0.06fF
C1387 greater comparator_0/NOR_0/w_0_0# 0.06fF
C1388 vdd addersubtractor_0/XOR_2/NAND_1/w_0_0# 0.05fF
C1389 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 gnd 0.11fF
C1390 twotofourdecoder_0/AND_3/NAND_0/a_6_n14# gnd 0.57fF
C1391 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_0_0# 0.05fF
C1392 twotofourdecoder_0/AND_2/not_0/w_0_0# vdd 0.05fF
C1393 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_0/a_6_n14# 0.12fF
C1394 addersubtractor_0/XOR_0/NAND_3/in1 addersubtractor_0/XOR_0/NAND_1/w_0_0# 0.03fF
C1395 enableblock_2/enable1_1/AND_1/NAND_0/a_6_n14# enableblock_2/enable1_1/AND_1/not_0/in 0.12fF
C1396 A0 enableblock_2/En 0.13fF
C1397 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_32_0# 0.05fF
C1398 gnd addersubtractor_0/fulladder_2/XOR_1/NAND_1/a_6_n14# 0.57fF
C1399 addersubtractor_0/XOR_0/NAND_3/w_32_0# addersubtractor_0/XOR_0/NAND_3/in2 0.06fF
C1400 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_32_0# addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 0.03fF
C1401 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_32_0# 0.05fF
C1402 addersubtractor_0/fulladder_2/XOR_0/NAND_1/a_6_n14# gnd 0.57fF
C1403 comparator_0/fourinputAND_1/fourinputNAND_0/w_100_0# comparator_0/XNOR_2/out 0.06fF
C1404 twotofourdecoder_0/AND_3/NAND_0/w_0_0# vdd 0.05fF
C1405 enableblock_2/enable1_0/AND_1/NAND_0/w_0_0# enableblock_2/enable1_0/AND_1/not_0/in 0.03fF
C1406 andblock_0/AND_3/not_0/in andblock_0/AND_3/NAND_0/w_0_0# 0.03fF
C1407 comparator_0/not_1/out comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# 0.02fF
C1408 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_0_0# 0.05fF
C1409 addersubtractor_0/XOR_2/out addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_32_0# 0.06fF
C1410 andblock_0/B2 gnd 0.38fF
C1411 andblock_0/A1 vdd 0.20fF
C1412 gnd addersubtractor_0/fulladder_3/XOR_1/in2 0.63fF
C1413 comparator_0/XNOR_0/XOR_0/NAND_1/w_0_0# comparator_0/XNOR_0/XOR_0/NAND_3/in1 0.03fF
C1414 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_0_0# 0.05fF
C1415 addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_32_0# addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 0.03fF
C1416 comparator_0/XNOR_1/XOR_0/NAND_3/w_0_0# comparator_0/XNOR_1/not_0/in 0.03fF
C1417 enableblock_2/enable1_0/AND_2/not_0/w_0_0# enableblock_2/enable1_0/AND_2/not_0/in 0.06fF
C1418 comparator_0/A2 comparator_0/B3 2.23fF
C1419 enableblock_1/enable1_0/AND_1/not_0/in enableblock_1/enable1_0/AND_1/NAND_0/a_6_n14# 0.12fF
C1420 addersubtractor_0/fulladder_0/OR_0/in2 vdd 0.07fF
C1421 vdd lesser 0.10fF
C1422 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_0/C 0.06fF
C1423 B0 enableblock_2/En 0.06fF
C1424 AND_2/not_0/w_0_0# AND_2/not_0/in 0.06fF
C1425 vdd addersubtractor_0/XOR_3/NAND_3/w_0_0# 0.05fF
C1426 comparator_0/XNOR_0/out comparator_0/fourinputAND_1/fourinputNAND_0/a_45_n14# 0.21fF
C1427 and0 gnd 0.08fF
C1428 enableblock_2/enable1_1/AND_0/NAND_0/a_6_n14# enableblock_2/enable1_1/AND_0/not_0/in 0.12fF
C1429 addersubtractor_0/fulladder_3/AND_0/not_0/in addersubtractor_0/fulladder_3/AND_0/NAND_0/a_6_n14# 0.12fF
C1430 comparator_0/not_2/out comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# 0.02fF
C1431 comparator_0/threeinputAND_0/not_0/w_0_0# vdd 0.05fF
C1432 comparator_0/fourinputAND_1/fourinputNAND_0/a_6_n14# gnd 0.47fF
C1433 andblock_0/AND_3/not_0/in vdd 0.29fF
C1434 comparator_0/XNOR_2/XOR_0/NAND_1/w_0_0# comparator_0/XNOR_2/XOR_0/NAND_3/in1 0.03fF
C1435 enableblock_1/enable1_0/AND_1/not_0/in gnd 0.04fF
C1436 addersubtractor_0/fulladder_3/AND_0/NAND_0/w_32_0# vdd 0.05fF
C1437 OR_0/NOT_0/in gnd 0.60fF
C1438 comparator_0/XNOR_0/XOR_0/NAND_3/w_0_0# comparator_0/XNOR_0/not_0/in 0.03fF
C1439 addersubtractor_0/XOR_3/NAND_2/w_32_0# addersubtractor_0/XOR_3/NAND_3/in2 0.03fF
C1440 OR_0/NOR_0/w_32_0# vdd 0.03fF
C1441 enableblock_0/A_out2 enableblock_0/enable1_0/AND_1/not_0/in 0.02fF
C1442 addersubtractor_0/XOR_1/out addersubtractor_0/XOR_1/NAND_3/w_0_0# 0.03fF
C1443 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_32_0# 0.03fF
C1444 comparator_0/XNOR_0/XOR_0/NAND_2/in1 gnd 0.15fF
C1445 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_0_0# vdd 0.05fF
C1446 comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# comparator_0/fourinputAND_0/fourinputNAND_0/a_45_n14# 0.04fF
C1447 comparator_0/fourinputAND_0/fourinputNAND_0/w_100_0# comparator_0/XNOR_0/out 0.06fF
C1448 enableblock_2/enable1_1/AND_3/NAND_0/w_32_0# enableblock_2/enable1_1/AND_3/not_0/in 0.03fF
C1449 and1 andblock_0/AND_2/not_0/in 0.02fF
C1450 andblock_0/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C1451 comparator_0/fourinputOR_0/in4 comparator_0/not_3/out 0.04fF
C1452 enableblock_0/enable1_1/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C1453 comparator_0/NOR_0/w_0_0# comparator_0/NOR_0/a_13_6# 0.03fF
C1454 comparator_0/XNOR_3/XOR_0/NAND_1/w_0_0# comparator_0/XNOR_3/XOR_0/NAND_3/in1 0.03fF
C1455 comparator_0/XNOR_1/XOR_0/NAND_0/w_32_0# comparator_0/XNOR_1/XOR_0/NAND_2/in1 0.03fF
C1456 gnd enableblock_1/enable1_0/AND_0/not_0/in 0.04fF
C1457 comparator_0/XNOR_2/XOR_0/NAND_3/w_0_0# comparator_0/XNOR_2/not_0/in 0.03fF
C1458 B1 AND_2/in2 0.06fF
C1459 addersubtractor_0/XOR_0/out addersubtractor_0/XOR_0/NAND_3/w_0_0# 0.03fF
C1460 OR_0/out OR_0/NOT_0/in 0.02fF
C1461 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_133_0# comparator_0/fiveinputAND_0/not_0/in 0.03fF
C1462 enableblock_1/enable1_1/AND_2/NAND_0/w_32_0# enableblock_1/enable1_1/AND_2/not_0/in 0.03fF
C1463 andblock_0/B2 andblock_0/AND_1/NAND_0/w_32_0# 0.06fF
C1464 comparator_0/NOR_0/w_32_0# comparator_0/NOR_0/a_13_6# 0.03fF
C1465 enableblock_0/enable1_0/AND_3/NAND_0/w_32_0# B1 0.06fF
C1466 comparator_0/fourinputAND_0/not_0/in gnd 0.01fF
C1467 enableblock_0/enable1_0/AND_0/not_0/in vdd 0.29fF
C1468 gnd addersubtractor_0/fulladder_3/AND_0/NAND_0/a_6_n14# 0.57fF
C1469 comparator_0/XNOR_1/XOR_0/NAND_3/in2 vdd 0.25fF
C1470 comparator_0/not_2/out vdd 0.07fF
C1471 comparator_0/fourinputAND_1/fourinputNAND_0/w_32_0# comparator_0/XNOR_0/out 0.06fF
C1472 addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_0/w_32_0# 0.03fF
C1473 comparator_0/XNOR_3/XOR_0/NAND_3/w_0_0# comparator_0/XNOR_3/not_0/in 0.03fF
C1474 comparator_0/XNOR_0/XOR_0/NAND_3/in2 vdd 0.25fF
C1475 comparator_0/threeinputAND_0/not_0/in gnd 0.75fF
C1476 andblock_0/B0 vdd 0.11fF
C1477 vdd addersubtractor_0/XOR_1/NAND_2/in1 0.25fF
C1478 addersubtractor_0/fulladder_3/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_3/AND_0/not_0/in 0.06fF
C1479 addersubtractor_0/fulladder_0/XOR_1/NAND_3/a_6_n14# gnd 0.57fF
C1480 enableblock_0/enable1_1/AND_2/not_0/in gnd 0.04fF
C1481 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_32_0# 0.05fF
C1482 comparator_0/XNOR_2/XOR_0/NAND_3/in2 vdd 0.25fF
C1483 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_76_n14# comparator_0/fiveinputAND_0/fiveinputNAND_0/a_113_n14# 0.04fF
C1484 comparator_0/not_2/w_0_0# comparator_0/B1 0.06fF
C1485 XOR_0/in1 vdd 0.07fF
C1486 B2 enableblock_2/enable1_0/AND_3/NAND_0/w_32_0# 0.06fF
C1487 B0 enableblock_2/enable1_1/AND_3/NAND_0/w_32_0# 0.06fF
C1488 addersubtractor_0/fulladder_0/XOR_0/NAND_3/a_6_n14# gnd 0.57fF
C1489 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_2/w_0_0# 0.06fF
C1490 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_32_0# vdd 0.05fF
C1491 XOR_0/NAND_0/w_0_0# XOR_0/in1 0.06fF
C1492 andblock_0/AND_1/not_0/in gnd 0.04fF
C1493 enableblock_0/A_out1 S0 0.06fF
C1494 comparator_0/XNOR_0/XOR_0/NAND_1/w_32_0# vdd 0.05fF
C1495 comparator_0/XNOR_0/out vdd 0.37fF
C1496 comparator_0/XNOR_1/XOR_0/NAND_1/w_32_0# comparator_0/XNOR_1/XOR_0/NAND_3/in1 0.03fF
C1497 enableblock_2/enable1_0/AND_1/not_0/w_0_0# andblock_0/B3 0.03fF
C1498 enableblock_0/enable1_1/AND_2/NAND_0/w_32_0# OR_0/out 0.06fF
C1499 addersubtractor_0/XOR_0/NAND_2/w_32_0# S0 0.06fF
C1500 comparator_0/XNOR_3/XOR_0/NAND_3/in2 vdd 0.25fF
C1501 enableblock_1/enable1_0/AND_3/NAND_0/w_32_0# enableblock_1/enable1_0/AND_3/not_0/in 0.03fF
C1502 AND_1/NAND_0/w_32_0# AND_1/in2 0.06fF
C1503 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 gnd 0.15fF
C1504 enableblock_0/enable1_0/AND_0/not_0/w_0_0# vdd 0.05fF
C1505 gnd addersubtractor_0/XOR_1/NAND_3/in1 0.11fF
C1506 comparator_0/XNOR_2/XOR_0/NAND_2/in1 gnd 0.15fF
C1507 addersubtractor_0/fulladder_1/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C1508 comparator_0/XNOR_2/XOR_0/NAND_1/w_32_0# vdd 0.05fF
C1509 gnd AND_0/in1 0.08fF
C1510 addersubtractor_0/fulladder_1/XOR_1/NAND_0/a_6_n14# gnd 0.57fF
C1511 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_32_0# addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 0.03fF
C1512 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_32_0# vdd 0.05fF
C1513 comparator_0/XNOR_1/XOR_0/NAND_2/w_0_0# comparator_0/XNOR_1/XOR_0/NAND_3/in2 0.03fF
C1514 vdd addersubtractor_0/fulladder_3/AND_1/not_0/in 0.29fF
C1515 addersubtractor_0/XOR_0/out gnd 0.56fF
C1516 comparator_0/A3 enableblock_1/enable1_0/AND_0/not_0/in 0.02fF
C1517 enableblock_0/B_out1 addersubtractor_0/XOR_3/out 0.11fF
C1518 vdd AND_0/not_0/w_0_0# 0.05fF
C1519 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_0_0# adder2 0.03fF
C1520 addersubtractor_0/fulladder_0/AND_0/NAND_0/w_32_0# vdd 0.05fF
C1521 addersubtractor_0/fulladder_0/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C1522 addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_0_0# 0.06fF
C1523 comparator_0/XNOR_3/XOR_0/NAND_1/w_32_0# vdd 0.05fF
C1524 comparator_0/XNOR_1/XOR_0/NAND_0/w_32_0# vdd 0.05fF
C1525 A2 B3 4.40fF
C1526 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 0.25fF
C1527 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_0_0# enableblock_0/A_out3 0.06fF
C1528 enableblock_2/enable1_0/AND_0/not_0/w_0_0# enableblock_2/enable1_0/AND_0/not_0/in 0.06fF
C1529 A0 B0 0.15fF
C1530 andblock_0/AND_2/NAND_0/a_6_n14# gnd 0.57fF
C1531 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_0/w_0_0# 0.03fF
C1532 vdd addersubtractor_0/fulladder_3/OR_0/NOR_0/w_0_0# 0.05fF
C1533 vdd addersubtractor_0/fulladder_0/C 0.18fF
C1534 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 0.25fF
C1535 S1 twotofourdecoder_0/not_1/out 0.16fF
C1536 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_0_0# addersubtractor_0/fulladder_2/XOR_1/in2 0.03fF
C1537 comparator_0/XNOR_0/XOR_0/NAND_2/w_0_0# comparator_0/XNOR_0/XOR_0/NAND_3/in2 0.03fF
C1538 enableblock_0/enable1_0/AND_1/NAND_0/w_0_0# vdd 0.05fF
C1539 vdd AND_0/NAND_0/w_32_0# 0.05fF
C1540 comparator_0/fourinputAND_0/not_0/w_0_0# vdd 0.05fF
C1541 comparator_0/not_0/out vdd 0.07fF
C1542 enableblock_2/enable1_1/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C1543 enableblock_0/enable1_0/AND_3/not_0/w_0_0# vdd 0.05fF
C1544 enableblock_0/enable1_1/AND_0/NAND_0/w_0_0# vdd 0.05fF
C1545 andblock_0/A0 enableblock_2/enable1_1/AND_2/not_0/in 0.02fF
C1546 A1 enableblock_2/enable1_1/AND_0/NAND_0/w_0_0# 0.06fF
C1547 enableblock_0/enable1_1/AND_0/not_0/in enableblock_0/enable1_1/AND_0/NAND_0/w_0_0# 0.03fF
C1548 addersubtractor_0/fulladder_1/XOR_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 0.12fF
C1549 addersubtractor_0/XOR_2/NAND_3/in1 addersubtractor_0/XOR_2/NAND_1/w_0_0# 0.03fF
C1550 andblock_0/AND_1/not_0/in andblock_0/AND_1/NAND_0/w_32_0# 0.03fF
C1551 comparator_0/A3 enableblock_1/enable1_0/AND_0/not_0/w_0_0# 0.03fF
C1552 comparator_0/XNOR_2/XOR_0/NAND_2/w_0_0# comparator_0/XNOR_2/XOR_0/NAND_3/in2 0.03fF
C1553 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 0.25fF
C1554 enableblock_0/enable1_0/AND_2/NAND_0/w_0_0# enableblock_0/enable1_0/AND_2/not_0/in 0.03fF
C1555 comparator_0/XNOR_1/XOR_0/NAND_2/a_6_n14# gnd 0.59fF
C1556 comparator_0/XNOR_1/XOR_0/NAND_2/w_32_0# vdd 0.05fF
C1557 enableblock_2/enable1_1/AND_2/NAND_0/a_6_n14# gnd 0.57fF
C1558 enableblock_2/enable1_1/AND_1/not_0/w_0_0# vdd 0.05fF
C1559 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_45_n14# comparator_0/A0 0.14fF
C1560 B3 enableblock_1/enable1_0/AND_1/NAND_0/w_32_0# 0.06fF
C1561 addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_32_0# 0.06fF
C1562 enableblock_0/enable1_0/AND_0/NAND_0/w_32_0# enableblock_0/enable1_0/AND_0/not_0/in 0.03fF
C1563 addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_32_0# 0.06fF
C1564 enableblock_0/enable1_0/AND_3/not_0/w_0_0# enableblock_0/enable1_0/AND_3/not_0/in 0.06fF
C1565 gnd enableblock_1/enable1_1/AND_1/NAND_0/a_6_n14# 0.57fF
C1566 S0 addersubtractor_0/XOR_3/NAND_0/w_32_0# 0.06fF
C1567 comparator_0/XNOR_3/XOR_0/NAND_2/w_0_0# comparator_0/XNOR_3/XOR_0/NAND_3/in2 0.03fF
C1568 comparator_0/XNOR_0/XOR_0/NAND_2/w_32_0# vdd 0.05fF
C1569 comparator_0/XNOR_0/XOR_0/NAND_2/a_6_n14# gnd 0.59fF
C1570 vdd enableblock_1/enable1_1/AND_0/not_0/w_0_0# 0.05fF
C1571 addersubtractor_0/fulladder_2/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C1572 vdd addersubtractor_0/fulladder_1/OR_0/in2 0.07fF
C1573 enableblock_2/enable1_1/AND_2/NAND_0/w_0_0# vdd 0.05fF
C1574 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_1/a_6_n14# 0.12fF
C1575 twotofourdecoder_0/AND_0/not_0/in gnd 0.04fF
C1576 enableblock_2/enable1_1/AND_3/NAND_0/w_0_0# enableblock_2/En 0.06fF
C1577 comparator_0/XNOR_2/XOR_0/NAND_2/w_32_0# vdd 0.05fF
C1578 comparator_0/XNOR_2/XOR_0/NAND_2/a_6_n14# gnd 0.59fF
C1579 B2 gnd 0.83fF
C1580 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_0_0# S0 0.06fF
C1581 and3 andblock_0/AND_0/not_0/in 0.02fF
C1582 vdd enableblock_1/enable1_1/AND_1/NAND_0/w_0_0# 0.05fF
C1583 addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_0/OR_0/NOR_0/w_32_0# 0.03fF
C1584 addersubtractor_0/fulladder_1/AND_1/not_0/in gnd 0.04fF
C1585 comparator_0/XNOR_3/XOR_0/NAND_2/a_6_n14# gnd 0.59fF
C1586 twotofourdecoder_0/AND_1/not_0/in gnd 0.04fF
C1587 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_1/a_6_n14# 0.12fF
C1588 comparator_0/XNOR_3/XOR_0/NAND_2/w_32_0# vdd 0.05fF
C1589 enableblock_0/B_out0 gnd 0.82fF
C1590 addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/OR_0/NOT_0/in 0.26fF
C1591 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_32_0# addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 0.03fF
C1592 vdd enableblock_1/enable1_1/AND_3/not_0/w_0_0# 0.05fF
C1593 enableblock_1/enable1_1/AND_1/NAND_0/w_0_0# AND_2/in2 0.06fF
C1594 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_0_0# 0.05fF
C1595 comparator_0/AND_0/NAND_0/w_32_0# vdd 0.05fF
C1596 addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_32_0# addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 0.03fF
C1597 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_0_0# 0.05fF
C1598 B2 OR_0/out 0.06fF
C1599 vdd enableblock_0/A_out1 0.32fF
C1600 enableblock_0/B_out1 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_0_0# 0.06fF
C1601 vdd addersubtractor_0/XOR_0/NAND_2/w_32_0# 0.05fF
C1602 enableblock_2/En twotofourdecoder_0/not_1/out 0.06fF
C1603 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_0_0# addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 0.03fF
C1604 gnd addersubtractor_0/fulladder_2/XOR_1/NAND_2/a_6_n14# 0.59fF
C1605 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_32_0# addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 0.03fF
C1606 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_32_0# 0.05fF
C1607 comparator_0/fourinputOR_0/in2 comparator_0/XNOR_1/out 0.06fF
C1608 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_32_0# 0.05fF
C1609 enableblock_2/enable1_0/AND_2/NAND_0/w_32_0# vdd 0.05fF
C1610 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_32_0# addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 0.06fF
C1611 vdd addersubtractor_0/fulladder_3/OR_0/NOT_0/in 0.11fF
C1612 addersubtractor_0/fulladder_3/OR_0/NOT_0/in addersubtractor_0/fulladder_3/OR_0/NOT_0/w_0_0# 0.06fF
C1613 addersubtractor_0/fulladder_2/XOR_0/NAND_2/a_6_n14# gnd 0.59fF
C1614 vdd addersubtractor_0/fulladder_1/OR_0/in1 0.12fF
C1615 comparator_0/AND_0/NAND_0/a_6_n14# comparator_0/AND_0/not_0/in 0.12fF
C1616 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_32_0# 0.05fF
C1617 enableblock_2/enable1_1/AND_1/not_0/w_0_0# enableblock_2/enable1_1/AND_1/not_0/in 0.06fF
C1618 addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_0_0# addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 0.03fF
C1619 OR_0/in1 XOR_0/NAND_2/w_32_0# 0.06fF
C1620 OR_0/in1 vdd 0.31fF
C1621 addersubtractor_0/fulladder_0/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_0/OR_0/in2 0.03fF
C1622 B3 A1 0.19fF
C1623 A3 B1 0.19fF
C1624 S1 gnd 0.78fF
C1625 enableblock_2/enable1_0/AND_2/not_0/in vdd 0.29fF
C1626 adder3 addersubtractor_0/fulladder_3/XOR_1/NAND_3/a_6_n14# 0.12fF
C1627 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 0.06fF
C1628 vdd AND_2/not_0/in 0.29fF
C1629 addersubtractor_0/fulladder_2/OR_0/NOT_0/in addersubtractor_0/fulladder_2/C 0.02fF
C1630 OR_0/in1 AND_2/in2 0.13fF
C1631 XOR_0/NAND_3/w_0_0# Carry 0.03fF
C1632 enableblock_1/enable1_1/AND_0/not_0/w_0_0# enableblock_1/enable1_1/AND_0/not_0/in 0.06fF
C1633 comparator_0/XNOR_2/out comparator_0/XNOR_2/not_0/w_0_0# 0.03fF
C1634 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_3/a_6_n14# 0.12fF
C1635 and1 vdd 0.20fF
C1636 gnd addersubtractor_0/XOR_3/NAND_1/a_6_n14# 0.57fF
C1637 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_0_0# 0.06fF
C1638 AND_2/NAND_0/a_6_n14# AND_2/not_0/in 0.12fF
C1639 vdd addersubtractor_0/XOR_3/NAND_1/w_32_0# 0.05fF
C1640 andblock_0/AND_2/NAND_0/a_6_n14# andblock_0/AND_2/not_0/in 0.12fF
C1641 comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_32_0# 0.03fF
C1642 addersubtractor_0/XOR_3/NAND_3/w_32_0# addersubtractor_0/XOR_3/NAND_3/in2 0.06fF
C1643 comparator_0/XNOR_0/XOR_0/NAND_1/w_32_0# comparator_0/XNOR_0/XOR_0/NAND_3/in1 0.03fF
C1644 enableblock_2/enable1_1/AND_1/NAND_0/w_32_0# vdd 0.05fF
C1645 enableblock_2/enable1_1/AND_3/NAND_0/w_0_0# enableblock_2/enable1_1/AND_3/not_0/in 0.03fF
C1646 XOR_0/NAND_3/in1 gnd 0.11fF
C1647 XOR_0/in1 AND_0/not_0/in 0.02fF
C1648 comparator_0/B1 enableblock_1/enable1_1/AND_1/not_0/w_0_0# 0.03fF
C1649 gnd addersubtractor_0/XOR_1/NAND_3/a_6_n14# 0.57fF
C1650 vdd addersubtractor_0/XOR_1/NAND_3/w_32_0# 0.05fF
C1651 enableblock_1/enable1_0/AND_1/not_0/w_0_0# enableblock_1/enable1_0/AND_1/not_0/in 0.06fF
C1652 enableblock_1/enable1_1/AND_2/NAND_0/w_0_0# enableblock_1/enable1_1/AND_2/not_0/in 0.03fF
C1653 XOR_0/NAND_1/w_0_0# vdd 0.05fF
C1654 comparator_0/B1 comparator_0/XNOR_1/out 0.07fF
C1655 comparator_0/XNOR_2/XOR_0/NAND_1/w_32_0# comparator_0/XNOR_2/XOR_0/NAND_3/in1 0.03fF
C1656 vdd addersubtractor_0/XOR_3/NAND_0/w_32_0# 0.05fF
C1657 andblock_0/AND_1/not_0/w_0_0# and2 0.03fF
C1658 comparator_0/fourinputAND_1/fourinputNAND_0/a_6_n14# comparator_0/fourinputAND_1/fourinputNAND_0/a_45_n14# 0.04fF
C1659 enableblock_1/enable1_1/AND_3/not_0/w_0_0# enableblock_1/enable1_1/AND_3/not_0/in 0.06fF
C1660 addersubtractor_0/fulladder_1/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_1/OR_0/in1 0.03fF
C1661 comparator_0/B0 comparator_0/XNOR_1/out 0.07fF
C1662 A0 enableblock_1/enable1_1/AND_2/NAND_0/w_0_0# 0.06fF
C1663 AND_0/not_0/in AND_0/not_0/w_0_0# 0.06fF
C1664 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_0_0# enableblock_0/A_out1 0.06fF
C1665 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_32_0# 0.06fF
C1666 addersubtractor_0/fulladder_2/AND_0/NAND_0/a_6_n14# addersubtractor_0/XOR_2/out 0.07fF
C1667 enableblock_0/B_out0 enableblock_0/enable1_1/AND_3/not_0/in 0.02fF
C1668 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_0_0# vdd 0.05fF
C1669 addersubtractor_0/fulladder_1/OR_0/NOT_0/in gnd 0.60fF
C1670 addersubtractor_0/fulladder_0/OR_0/NOT_0/in addersubtractor_0/fulladder_0/C 0.02fF
C1671 comparator_0/XNOR_3/XOR_0/NAND_1/w_32_0# comparator_0/XNOR_3/XOR_0/NAND_3/in1 0.03fF
C1672 OR_0/in2 gnd 0.34fF
C1673 addersubtractor_0/fulladder_3/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_2/C 0.07fF
C1674 addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_0_0# addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 0.03fF
C1675 enableblock_2/enable1_0/AND_0/NAND_0/w_32_0# enableblock_2/En 0.06fF
C1676 AND_0/not_0/in AND_0/NAND_0/w_32_0# 0.03fF
C1677 and2 vdd 0.18fF
C1678 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 0.25fF
C1679 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_0/w_32_0# 0.03fF
C1680 enableblock_2/En gnd 3.63fF
C1681 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_0_0# addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 0.03fF
C1682 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 0.25fF
C1683 AND_2/in1 comparator_0/NOR_0/w_32_0# 0.06fF
C1684 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_0/a_6_n14# 0.12fF
C1685 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_0_0# 0.06fF
C1686 vdd addersubtractor_0/fulladder_3/AND_1/NAND_0/w_0_0# 0.05fF
C1687 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_0_0# addersubtractor_0/fulladder_0/C 0.06fF
C1688 enableblock_2/enable1_1/AND_1/NAND_0/w_32_0# enableblock_2/enable1_1/AND_1/not_0/in 0.03fF
C1689 enableblock_1/enable1_0/AND_3/NAND_0/w_0_0# enableblock_1/enable1_0/AND_3/not_0/in 0.03fF
C1690 comparator_0/not_3/w_0_0# vdd 0.05fF
C1691 OR_0/out OR_0/in2 0.76fF
C1692 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_32_0# 0.06fF
C1693 comparator_0/fourinputOR_0/in2 comparator_0/XNOR_2/out 0.13fF
C1694 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_0_0# comparator_0/not_3/out 0.06fF
C1695 addersubtractor_0/fulladder_3/XOR_1/NAND_2/a_6_n14# addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 0.12fF
C1696 OR_0/NOR_0/a_13_6# OR_0/NOR_0/w_32_0# 0.03fF
C1697 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_32_0# vdd 0.05fF
C1698 addersubtractor_0/fulladder_0/AND_0/not_0/in gnd 0.04fF
C1699 XOR_0/NAND_2/w_0_0# XOR_0/NAND_3/in2 0.03fF
C1700 vdd adder3 0.25fF
C1701 andblock_0/AND_3/not_0/in andblock_0/AND_3/NAND_0/a_6_n14# 0.12fF
C1702 comparator_0/fourinputAND_1/fourinputNAND_0/w_0_0# comparator_0/XNOR_3/out 0.06fF
C1703 andblock_0/B2 vdd 0.17fF
C1704 addersubtractor_0/XOR_3/out addersubtractor_0/XOR_3/NAND_3/w_0_0# 0.03fF
C1705 vdd addersubtractor_0/fulladder_3/XOR_1/in2 0.47fF
C1706 addersubtractor_0/fulladder_3/XOR_0/NAND_2/a_6_n14# addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 0.12fF
C1707 comparator_0/fourinputOR_0/in2 gnd 0.16fF
C1708 comparator_0/XNOR_0/out comparator_0/B2 0.07fF
C1709 comparator_0/fourinputAND_0/fourinputNAND_0/w_100_0# comparator_0/fourinputAND_0/not_0/in 0.03fF
C1710 enableblock_0/enable1_0/AND_2/not_0/in gnd 0.04fF
C1711 comparator_0/fourinputAND_1/fourinputNAND_0/w_100_0# vdd 0.05fF
C1712 enableblock_1/enable1_0/AND_0/NAND_0/w_0_0# enableblock_1/enable1_0/AND_0/not_0/in 0.03fF
C1713 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_32_0# addersubtractor_0/XOR_0/out 0.06fF
C1714 OR_0/out enableblock_0/enable1_0/AND_2/NAND_0/w_32_0# 0.06fF
C1715 comparator_0/A2 gnd 1.18fF
C1716 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 0.15fF
C1717 and0 vdd 0.10fF
C1718 enableblock_2/enable1_1/AND_3/not_0/w_0_0# andblock_0/B0 0.03fF
C1719 comparator_0/XNOR_3/XOR_0/NAND_2/in1 gnd 0.15fF
C1720 comparator_0/fourinputAND_0/not_0/in comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# 0.11fF
C1721 enableblock_1/enable1_0/AND_1/not_0/in vdd 0.29fF
C1722 addersubtractor_0/XOR_3/NAND_2/a_6_n14# addersubtractor_0/XOR_3/NAND_3/in2 0.12fF
C1723 OR_0/NOT_0/in vdd 0.11fF
C1724 comparator_0/XNOR_1/XOR_0/NAND_0/w_32_0# comparator_0/B2 0.06fF
C1725 comparator_0/XNOR_0/XOR_0/NAND_2/in1 vdd 0.25fF
C1726 comparator_0/AND_0/not_0/w_0_0# comparator_0/AND_0/out 0.03fF
C1727 enableblock_0/enable1_1/AND_1/NAND_0/w_0_0# enableblock_0/enable1_1/AND_1/not_0/in 0.03fF
C1728 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_133_0# comparator_0/XNOR_2/out 0.06fF
C1729 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_63_0# comparator_0/fiveinputAND_0/not_0/in 0.03fF
C1730 A2 B1 0.23fF
C1731 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_32_0# adder0 0.03fF
C1732 enableblock_0/enable1_1/AND_2/not_0/w_0_0# enableblock_0/enable1_1/AND_2/not_0/in 0.06fF
C1733 comparator_0/XNOR_1/XOR_0/NAND_3/w_32_0# vdd 0.05fF
C1734 comparator_0/XNOR_1/XOR_0/NAND_3/a_6_n14# gnd 0.57fF
C1735 comparator_0/fourinputAND_0/fourinputNAND_0/w_63_0# vdd 0.05fF
C1736 vdd enableblock_1/enable1_0/AND_0/not_0/in 0.29fF
C1737 addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_0/w_0_0# 0.03fF
C1738 comparator_0/XNOR_2/out comparator_0/fiveinputAND_0/not_0/in 0.16fF
C1739 comparator_0/threeinputAND_0/threeinputNAND_0/a_45_n14# comparator_0/A2 0.18fF
C1740 comparator_0/XNOR_2/out comparator_0/B1 0.84fF
C1741 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_0/a_6_n14# 0.12fF
C1742 comparator_0/XNOR_0/XOR_0/NAND_3/a_6_n14# gnd 0.57fF
C1743 comparator_0/fourinputOR_0/fourinputNOR_0/w_32_0# comparator_0/fourinputOR_0/in2 0.06fF
C1744 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_0/XOR_1/in2 0.03fF
C1745 comparator_0/XNOR_0/XOR_0/NAND_3/w_32_0# vdd 0.05fF
C1746 comparator_0/XNOR_1/not_0/w_0_0# comparator_0/XNOR_1/not_0/in 0.06fF
C1747 enableblock_2/enable1_1/AND_3/not_0/in gnd 0.04fF
C1748 enableblock_0/enable1_0/AND_1/NAND_0/w_32_0# B0 0.06fF
C1749 enableblock_0/enable1_0/AND_0/NAND_0/w_0_0# A0 0.06fF
C1750 comparator_0/B3 gnd 0.35fF
C1751 comparator_0/fourinputAND_0/not_0/in vdd 1.27fF
C1752 enableblock_0/enable1_0/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C1753 A3 enableblock_1/enable1_0/AND_0/NAND_0/a_6_n14# 0.07fF
C1754 B2 S0 0.20fF
C1755 XOR_0/NAND_0/w_32_0# vdd 0.05fF
C1756 comparator_0/XNOR_2/out comparator_0/B0 0.06fF
C1757 comparator_0/XNOR_2/XOR_0/NAND_3/a_6_n14# gnd 0.57fF
C1758 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_45_n14# comparator_0/fiveinputAND_0/fiveinputNAND_0/a_76_n14# 0.04fF
C1759 andblock_0/AND_1/not_0/w_0_0# andblock_0/AND_1/not_0/in 0.06fF
C1760 comparator_0/XNOR_2/XOR_0/NAND_3/w_32_0# vdd 0.05fF
C1761 comparator_0/fiveinputAND_0/not_0/in gnd 0.01fF
C1762 enableblock_0/enable1_1/AND_2/NAND_0/w_32_0# vdd 0.05fF
C1763 gnd enableblock_1/enable1_1/AND_2/not_0/in 0.04fF
C1764 enableblock_1/enable1_0/AND_2/not_0/in comparator_0/A2 0.02fF
C1765 comparator_0/B1 gnd 0.23fF
C1766 andblock_0/AND_1/NAND_0/w_0_0# andblock_0/AND_1/not_0/in 0.03fF
C1767 addersubtractor_0/fulladder_3/AND_0/NAND_0/w_0_0# addersubtractor_0/fulladder_3/AND_0/not_0/in 0.03fF
C1768 andblock_0/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C1769 comparator_0/XNOR_3/XOR_0/NAND_3/w_32_0# vdd 0.05fF
C1770 comparator_0/XNOR_3/XOR_0/NAND_3/a_6_n14# gnd 0.57fF
C1771 comparator_0/B2 comparator_0/XNOR_1/XOR_0/NAND_2/w_32_0# 0.06fF
C1772 comparator_0/threeinputAND_0/not_0/in vdd 1.58fF
C1773 enableblock_0/B_out0 S0 0.06fF
C1774 enableblock_0/enable1_1/AND_2/not_0/in vdd 0.29fF
C1775 A0 gnd 0.23fF
C1776 twotofourdecoder_0/AND_3/NAND_0/w_32_0# twotofourdecoder_0/AND_3/not_0/in 0.03fF
C1777 comparator_0/B0 gnd 0.22fF
C1778 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_0_0# 0.05fF
C1779 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_1/AND_1/not_0/in 0.03fF
C1780 vdd enableblock_1/enable1_0/AND_0/not_0/w_0_0# 0.05fF
C1781 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_2/w_0_0# 0.06fF
C1782 addersubtractor_0/fulladder_1/XOR_1/in2 gnd 0.63fF
C1783 enableblock_2/enable1_0/AND_2/NAND_0/a_6_n14# gnd 0.57fF
C1784 enableblock_2/enable1_0/AND_1/not_0/w_0_0# vdd 0.05fF
C1785 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_0_0# 0.05fF
C1786 enableblock_0/A_out3 gnd 1.67fF
C1787 andblock_0/AND_1/not_0/in vdd 0.29fF
C1788 comparator_0/XNOR_1/XOR_0/NAND_3/in1 comparator_0/XNOR_1/XOR_0/NAND_1/a_6_n14# 0.12fF
C1789 comparator_0/fourinputOR_0/in4 comparator_0/fiveinputAND_0/not_0/w_0_0# 0.03fF
C1790 comparator_0/fourinputOR_0/in4 comparator_0/fourinputOR_0/not_0/in 0.10fF
C1791 comparator_0/fourinputAND_1/fourinputNAND_0/w_0_0# vdd 0.05fF
C1792 enableblock_0/enable1_0/AND_2/not_0/w_0_0# enableblock_0/A_out1 0.03fF
C1793 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 0.25fF
C1794 XOR_0/NAND_2/w_0_0# vdd 0.05fF
C1795 vdd addersubtractor_0/XOR_1/NAND_3/in1 0.25fF
C1796 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_32_0# 0.05fF
C1797 gnd addersubtractor_0/fulladder_2/XOR_1/NAND_3/a_6_n14# 0.57fF
C1798 vdd addersubtractor_0/XOR_0/out 0.06fF
C1799 comparator_0/XNOR_2/XOR_0/NAND_2/in1 vdd 0.25fF
C1800 addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_3/OR_0/NOR_0/w_0_0# 0.03fF
C1801 greater gnd 0.08fF
C1802 enableblock_2/enable1_0/AND_2/NAND_0/w_0_0# vdd 0.05fF
C1803 AND_0/in1 addersubtractor_0/fulladder_3/OR_0/NOT_0/w_0_0# 0.03fF
C1804 vdd AND_0/in1 0.10fF
C1805 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_32_0# 0.05fF
C1806 addersubtractor_0/fulladder_2/XOR_0/NAND_3/a_6_n14# gnd 0.57fF
C1807 enableblock_2/En enableblock_2/enable1_0/AND_3/NAND_0/w_0_0# 0.06fF
C1808 B0 gnd 0.76fF
C1809 addersubtractor_0/XOR_0/out vdd 0.32fF
C1810 gnd AND_1/not_0/in 0.04fF
C1811 comparator_0/fourinputOR_0/in3 gnd 0.79fF
C1812 vdd enableblock_1/enable1_0/AND_1/NAND_0/w_0_0# 0.05fF
C1813 vdd AND_2/NAND_0/w_32_0# 0.05fF
C1814 comparator_0/XNOR_0/XOR_0/NAND_3/in1 comparator_0/XNOR_0/XOR_0/NAND_1/a_6_n14# 0.12fF
C1815 AND_1/not_0/w_0_0# AND_1/not_0/in 0.06fF
C1816 enableblock_0/A_out0 gnd 0.82fF
C1817 addersubtractor_0/fulladder_3/OR_0/NOT_0/in addersubtractor_0/fulladder_3/OR_0/NOR_0/w_32_0# 0.03fF
C1818 addersubtractor_0/XOR_0/NAND_2/a_6_n14# gnd 0.59fF
C1819 comparator_0/A3 comparator_0/B3 0.38fF
C1820 AND_2/NAND_0/w_32_0# AND_2/in2 0.06fF
C1821 vdd addersubtractor_0/fulladder_3/AND_0/not_0/w_0_0# 0.05fF
C1822 enableblock_1/enable1_0/AND_1/NAND_0/w_0_0# AND_2/in2 0.06fF
C1823 OR_0/out B0 0.06fF
C1824 enableblock_0/enable1_1/AND_1/not_0/w_0_0# enableblock_0/B_out2 0.03fF
C1825 comparator_0/XNOR_2/XOR_0/NAND_3/in1 comparator_0/XNOR_2/XOR_0/NAND_1/a_6_n14# 0.12fF
C1826 gnd addersubtractor_0/XOR_3/NAND_3/in1 0.11fF
C1827 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_0_0# addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 0.03fF
C1828 addersubtractor_0/XOR_0/NAND_2/w_32_0# addersubtractor_0/XOR_0/NAND_3/in2 0.03fF
C1829 A2 enableblock_0/enable1_1/AND_0/NAND_0/w_0_0# 0.06fF
C1830 twotofourdecoder_0/AND_0/NAND_0/w_32_0# twotofourdecoder_0/AND_0/not_0/in 0.03fF
C1831 comparator_0/A1 comparator_0/B1 0.95fF
C1832 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_32_0# addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 0.03fF
C1833 enableblock_0/enable1_0/AND_2/NAND_0/a_6_n14# enableblock_0/enable1_0/AND_2/not_0/in 0.12fF
C1834 andblock_0/B1 gnd 0.38fF
C1835 comparator_0/A0 enableblock_1/enable1_1/AND_2/not_0/in 0.02fF
C1836 comparator_0/AND_0/out comparator_0/fourinputOR_0/in2 1.17fF
C1837 addersubtractor_0/fulladder_2/XOR_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 0.12fF
C1838 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_32_0# addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 0.03fF
C1839 A1 B1 0.23fF
C1840 comparator_0/XNOR_3/XOR_0/NAND_3/in1 comparator_0/XNOR_3/XOR_0/NAND_1/a_6_n14# 0.12fF
C1841 comparator_0/A0 comparator_0/B0 0.13fF
C1842 addersubtractor_0/fulladder_1/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_1/OR_0/in2 0.03fF
C1843 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_2/w_0_0# 0.06fF
C1844 OR_0/NOT_0/in Gnd 0.77fF
C1845 OR_0/NOR_0/a_13_6# Gnd 0.02fF
C1846 OR_0/NOR_0/w_32_0# Gnd 0.40fF
C1847 OR_0/NOR_0/w_0_0# Gnd 0.40fF
C1848 OR_0/NOT_0/w_0_0# Gnd 0.40fF
C1849 XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C1850 Carry Gnd 0.53fF
C1851 XOR_0/NAND_3/in2 Gnd 0.76fF
C1852 XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C1853 XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C1854 XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C1855 XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C1856 XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C1857 XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C1858 XOR_0/NAND_3/in1 Gnd 0.78fF
C1859 XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C1860 XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C1861 XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C1862 XOR_0/NAND_2/in1 Gnd 0.97fF
C1863 XOR_0/in1 Gnd 1.72fF
C1864 XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C1865 XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C1866 andblock_0/AND_3/not_0/in Gnd 0.76fF
C1867 and0 Gnd 0.19fF
C1868 andblock_0/AND_3/not_0/w_0_0# Gnd 0.40fF
C1869 andblock_0/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C1870 andblock_0/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C1871 andblock_0/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C1872 andblock_0/AND_2/not_0/in Gnd 0.76fF
C1873 and1 Gnd 0.20fF
C1874 andblock_0/AND_2/not_0/w_0_0# Gnd 0.40fF
C1875 andblock_0/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C1876 andblock_0/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C1877 andblock_0/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C1878 andblock_0/AND_1/not_0/in Gnd 0.76fF
C1879 and2 Gnd 0.20fF
C1880 andblock_0/AND_1/not_0/w_0_0# Gnd 0.40fF
C1881 andblock_0/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C1882 andblock_0/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C1883 andblock_0/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C1884 andblock_0/AND_0/not_0/in Gnd 0.76fF
C1885 and3 Gnd 0.20fF
C1886 andblock_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C1887 andblock_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C1888 andblock_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C1889 andblock_0/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C1890 comparator_0/NOR_0/a_13_6# Gnd 0.02fF
C1891 comparator_0/NOR_0/w_32_0# Gnd 0.40fF
C1892 comparator_0/NOR_0/w_0_0# Gnd 0.40fF
C1893 comparator_0/XNOR_3/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C1894 comparator_0/XNOR_3/not_0/in Gnd 0.76fF
C1895 comparator_0/XNOR_3/XOR_0/NAND_3/in2 Gnd 0.76fF
C1896 comparator_0/XNOR_3/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C1897 comparator_0/XNOR_3/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C1898 comparator_0/XNOR_3/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C1899 comparator_0/XNOR_3/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C1900 comparator_0/XNOR_3/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C1901 comparator_0/XNOR_3/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C1902 comparator_0/XNOR_3/XOR_0/NAND_3/in1 Gnd 0.78fF
C1903 comparator_0/XNOR_3/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C1904 comparator_0/XNOR_3/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C1905 comparator_0/XNOR_3/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C1906 comparator_0/XNOR_3/XOR_0/NAND_2/in1 Gnd 0.97fF
C1907 comparator_0/B0 Gnd 1.82fF
C1908 comparator_0/A0 Gnd 3.08fF
C1909 comparator_0/XNOR_3/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C1910 comparator_0/XNOR_3/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C1911 comparator_0/XNOR_3/not_0/w_0_0# Gnd 0.40fF
C1912 comparator_0/XNOR_2/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C1913 comparator_0/XNOR_2/not_0/in Gnd 0.76fF
C1914 comparator_0/XNOR_2/XOR_0/NAND_3/in2 Gnd 0.76fF
C1915 comparator_0/XNOR_2/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C1916 comparator_0/XNOR_2/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C1917 comparator_0/XNOR_2/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C1918 comparator_0/XNOR_2/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C1919 comparator_0/XNOR_2/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C1920 comparator_0/XNOR_2/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C1921 comparator_0/XNOR_2/XOR_0/NAND_3/in1 Gnd 0.78fF
C1922 comparator_0/XNOR_2/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C1923 comparator_0/XNOR_2/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C1924 comparator_0/XNOR_2/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C1925 comparator_0/XNOR_2/XOR_0/NAND_2/in1 Gnd 0.97fF
C1926 comparator_0/B1 Gnd 1.62fF
C1927 comparator_0/A1 Gnd 2.60fF
C1928 comparator_0/XNOR_2/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C1929 comparator_0/XNOR_2/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C1930 comparator_0/XNOR_2/not_0/w_0_0# Gnd 0.40fF
C1931 comparator_0/XNOR_0/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C1932 comparator_0/XNOR_0/not_0/in Gnd 0.76fF
C1933 comparator_0/XNOR_0/XOR_0/NAND_3/in2 Gnd 0.76fF
C1934 comparator_0/XNOR_0/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C1935 comparator_0/XNOR_0/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C1936 comparator_0/XNOR_0/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C1937 comparator_0/XNOR_0/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C1938 comparator_0/XNOR_0/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C1939 comparator_0/XNOR_0/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C1940 comparator_0/XNOR_0/XOR_0/NAND_3/in1 Gnd 0.78fF
C1941 comparator_0/XNOR_0/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C1942 comparator_0/XNOR_0/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C1943 comparator_0/XNOR_0/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C1944 comparator_0/XNOR_0/XOR_0/NAND_2/in1 Gnd 0.97fF
C1945 comparator_0/B3 Gnd 0.01fF
C1946 comparator_0/A3 Gnd 1.29fF
C1947 comparator_0/XNOR_0/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C1948 comparator_0/XNOR_0/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C1949 comparator_0/XNOR_0/not_0/w_0_0# Gnd 0.40fF
C1950 comparator_0/XNOR_1/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C1951 comparator_0/XNOR_1/not_0/in Gnd 0.76fF
C1952 comparator_0/XNOR_1/XOR_0/NAND_3/in2 Gnd 0.76fF
C1953 comparator_0/XNOR_1/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C1954 comparator_0/XNOR_1/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C1955 comparator_0/XNOR_1/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C1956 comparator_0/XNOR_1/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C1957 comparator_0/XNOR_1/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C1958 comparator_0/XNOR_1/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C1959 comparator_0/XNOR_1/XOR_0/NAND_3/in1 Gnd 0.78fF
C1960 comparator_0/XNOR_1/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C1961 comparator_0/XNOR_1/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C1962 comparator_0/XNOR_1/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C1963 comparator_0/XNOR_1/XOR_0/NAND_2/in1 Gnd 0.97fF
C1964 comparator_0/B2 Gnd 2.68fF
C1965 comparator_0/A2 Gnd 2.23fF
C1966 comparator_0/XNOR_1/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C1967 comparator_0/XNOR_1/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C1968 comparator_0/XNOR_1/not_0/w_0_0# Gnd 0.40fF
C1969 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_113_n14# Gnd 0.08fF
C1970 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_76_n14# Gnd 0.05fF
C1971 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_45_n14# Gnd 0.07fF
C1972 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# Gnd 0.14fF
C1973 comparator_0/fiveinputAND_0/not_0/in Gnd 1.48fF
C1974 comparator_0/XNOR_2/out Gnd 1.52fF
C1975 comparator_0/not_3/out Gnd 1.44fF
C1976 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_133_0# Gnd 0.43fF
C1977 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_63_0# Gnd 0.43fF
C1978 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_32_0# Gnd 0.43fF
C1979 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_0_0# Gnd 0.43fF
C1980 comparator_0/fiveinputAND_0/not_0/w_0_0# Gnd 0.40fF
C1981 comparator_0/fourinputOR_0/in2 Gnd 1.03fF
C1982 comparator_0/threeinputAND_0/not_0/w_0_0# Gnd 0.40fF
C1983 comparator_0/threeinputAND_0/threeinputNAND_0/a_45_n14# Gnd 0.07fF
C1984 comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# Gnd 0.14fF
C1985 comparator_0/XNOR_0/out Gnd 0.53fF
C1986 comparator_0/not_1/out Gnd 0.29fF
C1987 comparator_0/threeinputAND_0/not_0/in Gnd 0.76fF
C1988 comparator_0/threeinputAND_0/threeinputNAND_0/w_63_0# Gnd 0.39fF
C1989 comparator_0/threeinputAND_0/threeinputNAND_0/w_32_0# Gnd 0.40fF
C1990 comparator_0/threeinputAND_0/threeinputNAND_0/w_0_0# Gnd 0.40fF
C1991 comparator_0/fourinputAND_1/fourinputNAND_0/a_76_n14# Gnd 0.05fF
C1992 comparator_0/fourinputAND_1/fourinputNAND_0/a_45_n14# Gnd 0.07fF
C1993 comparator_0/fourinputAND_1/fourinputNAND_0/a_6_n14# Gnd 0.14fF
C1994 comparator_0/fourinputAND_1/not_0/in Gnd 1.84fF
C1995 comparator_0/XNOR_3/out Gnd 0.61fF
C1996 comparator_0/fourinputAND_1/fourinputNAND_0/w_100_0# Gnd 0.40fF
C1997 comparator_0/fourinputAND_1/fourinputNAND_0/w_63_0# Gnd 0.40fF
C1998 comparator_0/fourinputAND_1/fourinputNAND_0/w_32_0# Gnd 0.40fF
C1999 comparator_0/fourinputAND_1/fourinputNAND_0/w_0_0# Gnd 0.40fF
C2000 comparator_0/fourinputAND_1/not_0/w_0_0# Gnd 0.40fF
C2001 comparator_0/fourinputAND_0/fourinputNAND_0/a_76_n14# Gnd 0.05fF
C2002 comparator_0/fourinputAND_0/fourinputNAND_0/a_45_n14# Gnd 0.07fF
C2003 comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# Gnd 0.14fF
C2004 comparator_0/fourinputAND_0/not_0/in Gnd 1.84fF
C2005 comparator_0/not_2/out Gnd 0.30fF
C2006 comparator_0/fourinputAND_0/fourinputNAND_0/w_100_0# Gnd 0.40fF
C2007 comparator_0/fourinputAND_0/fourinputNAND_0/w_63_0# Gnd 0.40fF
C2008 comparator_0/fourinputAND_0/fourinputNAND_0/w_32_0# Gnd 0.40fF
C2009 comparator_0/fourinputAND_0/fourinputNAND_0/w_0_0# Gnd 0.40fF
C2010 comparator_0/fourinputOR_0/in3 Gnd 1.03fF
C2011 comparator_0/fourinputAND_0/not_0/w_0_0# Gnd 0.40fF
C2012 comparator_0/not_3/w_0_0# Gnd 0.40fF
C2013 comparator_0/not_2/w_0_0# Gnd 0.40fF
C2014 comparator_0/not_1/w_0_0# Gnd 0.40fF
C2015 comparator_0/not_0/w_0_0# Gnd 0.40fF
C2016 comparator_0/AND_0/not_0/in Gnd 0.76fF
C2017 comparator_0/AND_0/out Gnd 1.01fF
C2018 comparator_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C2019 comparator_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2020 comparator_0/not_0/out Gnd 0.28fF
C2021 comparator_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2022 comparator_0/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2023 greater Gnd 1.58fF
C2024 comparator_0/fourinputOR_0/not_0/w_0_0# Gnd 0.40fF
C2025 comparator_0/fourinputOR_0/not_0/in Gnd 1.09fF
C2026 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# Gnd 0.02fF
C2027 comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# Gnd 0.02fF
C2028 comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# Gnd 0.02fF
C2029 comparator_0/fourinputOR_0/in4 Gnd 0.13fF
C2030 comparator_0/fourinputOR_0/fourinputNOR_0/w_97_0# Gnd 0.03fF
C2031 comparator_0/fourinputOR_0/fourinputNOR_0/w_64_0# Gnd 0.40fF
C2032 comparator_0/fourinputOR_0/fourinputNOR_0/w_32_0# Gnd 0.40fF
C2033 comparator_0/fourinputOR_0/fourinputNOR_0/w_0_0# Gnd 0.40fF
C2034 twotofourdecoder_0/not_1/w_0_0# Gnd 0.40fF
C2035 twotofourdecoder_0/not_0/w_0_0# Gnd 0.40fF
C2036 twotofourdecoder_0/AND_3/not_0/in Gnd 0.76fF
C2037 twotofourdecoder_0/AND_3/not_0/w_0_0# Gnd 0.40fF
C2038 twotofourdecoder_0/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2039 twotofourdecoder_0/not_1/out Gnd 1.39fF
C2040 twotofourdecoder_0/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2041 twotofourdecoder_0/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2042 twotofourdecoder_0/AND_2/not_0/in Gnd 0.76fF
C2043 OR_0/in2 Gnd 4.82fF
C2044 twotofourdecoder_0/AND_2/not_0/w_0_0# Gnd 0.40fF
C2045 twotofourdecoder_0/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2046 twotofourdecoder_0/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2047 twotofourdecoder_0/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2048 twotofourdecoder_0/AND_1/not_0/in Gnd 0.76fF
C2049 twotofourdecoder_0/AND_1/not_0/w_0_0# Gnd 0.40fF
C2050 twotofourdecoder_0/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2051 twotofourdecoder_0/not_0/out Gnd 1.67fF
C2052 twotofourdecoder_0/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2053 twotofourdecoder_0/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2054 twotofourdecoder_0/AND_0/not_0/in Gnd 0.76fF
C2055 twotofourdecoder_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C2056 twotofourdecoder_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2057 S1 Gnd 1.63fF
C2058 twotofourdecoder_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2059 twotofourdecoder_0/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2060 enableblock_2/enable1_0/AND_3/not_0/in Gnd 0.76fF
C2061 andblock_0/B2 Gnd 0.43fF
C2062 enableblock_2/enable1_0/AND_3/not_0/w_0_0# Gnd 0.40fF
C2063 enableblock_2/enable1_0/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2064 enableblock_2/enable1_0/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2065 enableblock_2/enable1_0/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2066 enableblock_2/enable1_0/AND_2/not_0/in Gnd 0.76fF
C2067 andblock_0/A2 Gnd 0.78fF
C2068 enableblock_2/enable1_0/AND_2/not_0/w_0_0# Gnd 0.40fF
C2069 enableblock_2/enable1_0/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2070 enableblock_2/enable1_0/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2071 enableblock_2/enable1_0/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2072 enableblock_2/enable1_0/AND_1/not_0/in Gnd 0.76fF
C2073 andblock_0/B3 Gnd 1.61fF
C2074 enableblock_2/enable1_0/AND_1/not_0/w_0_0# Gnd 0.40fF
C2075 enableblock_2/enable1_0/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2076 enableblock_2/En Gnd 5.01fF
C2077 enableblock_2/enable1_0/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2078 enableblock_2/enable1_0/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2079 enableblock_2/enable1_0/AND_0/not_0/in Gnd 0.76fF
C2080 enableblock_2/enable1_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C2081 enableblock_2/enable1_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2082 enableblock_2/enable1_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2083 enableblock_2/enable1_0/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2084 enableblock_2/enable1_1/AND_3/not_0/in Gnd 0.76fF
C2085 andblock_0/B0 Gnd 0.49fF
C2086 enableblock_2/enable1_1/AND_3/not_0/w_0_0# Gnd 0.40fF
C2087 enableblock_2/enable1_1/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2088 enableblock_2/enable1_1/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2089 enableblock_2/enable1_1/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2090 enableblock_2/enable1_1/AND_2/not_0/in Gnd 0.76fF
C2091 andblock_0/A0 Gnd 0.33fF
C2092 enableblock_2/enable1_1/AND_2/not_0/w_0_0# Gnd 0.40fF
C2093 enableblock_2/enable1_1/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2094 enableblock_2/enable1_1/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2095 enableblock_2/enable1_1/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2096 enableblock_2/enable1_1/AND_1/not_0/in Gnd 0.76fF
C2097 andblock_0/B1 Gnd 1.33fF
C2098 enableblock_2/enable1_1/AND_1/not_0/w_0_0# Gnd 0.40fF
C2099 enableblock_2/enable1_1/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2100 enableblock_2/enable1_1/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2101 enableblock_2/enable1_1/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2102 enableblock_2/enable1_1/AND_0/not_0/in Gnd 0.76fF
C2103 andblock_0/A1 Gnd 0.86fF
C2104 enableblock_2/enable1_1/AND_0/not_0/w_0_0# Gnd 0.40fF
C2105 enableblock_2/enable1_1/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2106 enableblock_2/enable1_1/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2107 enableblock_2/enable1_1/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2108 enableblock_0/enable1_0/AND_3/not_0/in Gnd 0.76fF
C2109 enableblock_0/A_out0 Gnd 1.45fF
C2110 enableblock_0/enable1_0/AND_3/not_0/w_0_0# Gnd 0.40fF
C2111 enableblock_0/enable1_0/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2112 B1 Gnd 40.05fF
C2113 enableblock_0/enable1_0/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2114 enableblock_0/enable1_0/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2115 enableblock_0/enable1_0/AND_2/not_0/in Gnd 0.76fF
C2116 enableblock_0/enable1_0/AND_2/not_0/w_0_0# Gnd 0.40fF
C2117 enableblock_0/enable1_0/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2118 A1 Gnd 1.13fF
C2119 enableblock_0/enable1_0/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2120 enableblock_0/enable1_0/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2121 enableblock_0/enable1_0/AND_1/not_0/in Gnd 0.76fF
C2122 enableblock_0/A_out2 Gnd 1.63fF
C2123 enableblock_0/enable1_0/AND_1/not_0/w_0_0# Gnd 0.40fF
C2124 enableblock_0/enable1_0/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2125 B0 Gnd 39.80fF
C2126 OR_0/out Gnd 5.23fF
C2127 enableblock_0/enable1_0/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2128 enableblock_0/enable1_0/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2129 enableblock_0/enable1_0/AND_0/not_0/in Gnd 0.76fF
C2130 enableblock_0/enable1_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C2131 enableblock_0/enable1_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2132 A0 Gnd 1.27fF
C2133 enableblock_0/enable1_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2134 enableblock_0/enable1_0/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2135 enableblock_0/enable1_1/AND_3/not_0/in Gnd 0.76fF
C2136 enableblock_0/B_out0 Gnd 0.22fF
C2137 enableblock_0/enable1_1/AND_3/not_0/w_0_0# Gnd 0.40fF
C2138 enableblock_0/enable1_1/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2139 B3 Gnd 40.94fF
C2140 enableblock_0/enable1_1/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2141 enableblock_0/enable1_1/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2142 enableblock_0/enable1_1/AND_2/not_0/in Gnd 0.76fF
C2143 enableblock_0/enable1_1/AND_2/not_0/w_0_0# Gnd 0.40fF
C2144 enableblock_0/enable1_1/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2145 A3 Gnd 1.15fF
C2146 enableblock_0/enable1_1/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2147 enableblock_0/enable1_1/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2148 enableblock_0/enable1_1/AND_1/not_0/in Gnd 0.76fF
C2149 enableblock_0/B_out2 Gnd 1.70fF
C2150 enableblock_0/enable1_1/AND_1/not_0/w_0_0# Gnd 0.40fF
C2151 enableblock_0/enable1_1/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2152 B2 Gnd 40.41fF
C2153 enableblock_0/enable1_1/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2154 enableblock_0/enable1_1/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2155 enableblock_0/enable1_1/AND_0/not_0/in Gnd 0.76fF
C2156 enableblock_0/enable1_1/AND_0/not_0/w_0_0# Gnd 0.40fF
C2157 enableblock_0/enable1_1/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2158 A2 Gnd 39.38fF
C2159 enableblock_0/enable1_1/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2160 enableblock_0/enable1_1/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2161 enableblock_1/enable1_0/AND_3/not_0/in Gnd 0.76fF
C2162 enableblock_1/enable1_0/AND_3/not_0/w_0_0# Gnd 0.40fF
C2163 enableblock_1/enable1_0/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2164 enableblock_1/enable1_0/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2165 enableblock_1/enable1_0/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2166 enableblock_1/enable1_0/AND_2/not_0/in Gnd 0.76fF
C2167 enableblock_1/enable1_0/AND_2/not_0/w_0_0# Gnd 0.40fF
C2168 enableblock_1/enable1_0/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2169 enableblock_1/enable1_0/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2170 enableblock_1/enable1_0/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2171 enableblock_1/enable1_0/AND_1/not_0/in Gnd 0.76fF
C2172 enableblock_1/enable1_0/AND_1/not_0/w_0_0# Gnd 0.40fF
C2173 enableblock_1/enable1_0/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2174 AND_2/in2 Gnd 15.07fF
C2175 enableblock_1/enable1_0/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2176 enableblock_1/enable1_0/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2177 enableblock_1/enable1_0/AND_0/not_0/in Gnd 0.76fF
C2178 enableblock_1/enable1_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C2179 enableblock_1/enable1_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2180 enableblock_1/enable1_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2181 enableblock_1/enable1_0/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2182 enableblock_1/enable1_1/AND_3/not_0/in Gnd 0.76fF
C2183 enableblock_1/enable1_1/AND_3/not_0/w_0_0# Gnd 0.40fF
C2184 enableblock_1/enable1_1/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2185 enableblock_1/enable1_1/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2186 enableblock_1/enable1_1/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2187 enableblock_1/enable1_1/AND_2/not_0/in Gnd 0.76fF
C2188 enableblock_1/enable1_1/AND_2/not_0/w_0_0# Gnd 0.40fF
C2189 enableblock_1/enable1_1/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2190 enableblock_1/enable1_1/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2191 enableblock_1/enable1_1/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2192 enableblock_1/enable1_1/AND_1/not_0/in Gnd 0.76fF
C2193 enableblock_1/enable1_1/AND_1/not_0/w_0_0# Gnd 0.40fF
C2194 enableblock_1/enable1_1/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2195 enableblock_1/enable1_1/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2196 enableblock_1/enable1_1/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2197 enableblock_1/enable1_1/AND_0/not_0/in Gnd 0.76fF
C2198 enableblock_1/enable1_1/AND_0/not_0/w_0_0# Gnd 0.40fF
C2199 enableblock_1/enable1_1/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2200 enableblock_1/enable1_1/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2201 enableblock_1/enable1_1/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2202 AND_2/not_0/in Gnd 0.76fF
C2203 equal Gnd 0.17fF
C2204 AND_2/not_0/w_0_0# Gnd 0.40fF
C2205 AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2206 AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2207 AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2208 AND_1/not_0/in Gnd 0.76fF
C2209 lesser Gnd 0.16fF
C2210 AND_1/not_0/w_0_0# Gnd 0.40fF
C2211 AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2212 AND_1/in2 Gnd 1.14fF
C2213 AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2214 AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2215 AND_0/not_0/in Gnd 0.76fF
C2216 AND_0/not_0/w_0_0# Gnd 0.40fF
C2217 AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2218 AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2219 AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2220 addersubtractor_0/XOR_3/NAND_3/a_6_n14# Gnd 0.14fF
C2221 addersubtractor_0/XOR_3/NAND_3/in2 Gnd 0.76fF
C2222 addersubtractor_0/XOR_3/NAND_3/w_32_0# Gnd 0.40fF
C2223 addersubtractor_0/XOR_3/NAND_3/w_0_0# Gnd 0.40fF
C2224 addersubtractor_0/XOR_3/NAND_2/a_6_n14# Gnd 0.14fF
C2225 addersubtractor_0/XOR_3/NAND_2/w_32_0# Gnd 0.40fF
C2226 addersubtractor_0/XOR_3/NAND_2/w_0_0# Gnd 0.40fF
C2227 addersubtractor_0/XOR_3/NAND_1/a_6_n14# Gnd 0.14fF
C2228 addersubtractor_0/XOR_3/NAND_3/in1 Gnd 0.78fF
C2229 addersubtractor_0/XOR_3/NAND_1/w_32_0# Gnd 0.40fF
C2230 addersubtractor_0/XOR_3/NAND_1/w_0_0# Gnd 0.40fF
C2231 addersubtractor_0/XOR_3/NAND_0/a_6_n14# Gnd 0.14fF
C2232 addersubtractor_0/XOR_3/NAND_2/in1 Gnd 0.97fF
C2233 addersubtractor_0/XOR_3/NAND_0/w_32_0# Gnd 0.40fF
C2234 addersubtractor_0/XOR_3/NAND_0/w_0_0# Gnd 0.40fF
C2235 addersubtractor_0/XOR_2/NAND_3/a_6_n14# Gnd 0.14fF
C2236 addersubtractor_0/XOR_2/NAND_3/in2 Gnd 0.76fF
C2237 addersubtractor_0/XOR_2/NAND_3/w_32_0# Gnd 0.40fF
C2238 addersubtractor_0/XOR_2/NAND_3/w_0_0# Gnd 0.40fF
C2239 addersubtractor_0/XOR_2/NAND_2/a_6_n14# Gnd 0.14fF
C2240 addersubtractor_0/XOR_2/NAND_2/w_32_0# Gnd 0.40fF
C2241 addersubtractor_0/XOR_2/NAND_2/w_0_0# Gnd 0.40fF
C2242 addersubtractor_0/XOR_2/NAND_1/a_6_n14# Gnd 0.14fF
C2243 addersubtractor_0/XOR_2/NAND_3/in1 Gnd 0.78fF
C2244 addersubtractor_0/XOR_2/NAND_1/w_32_0# Gnd 0.40fF
C2245 addersubtractor_0/XOR_2/NAND_1/w_0_0# Gnd 0.40fF
C2246 addersubtractor_0/XOR_2/NAND_0/a_6_n14# Gnd 0.14fF
C2247 addersubtractor_0/XOR_2/NAND_2/in1 Gnd 0.97fF
C2248 addersubtractor_0/XOR_2/NAND_0/w_32_0# Gnd 0.40fF
C2249 addersubtractor_0/XOR_2/NAND_0/w_0_0# Gnd 0.40fF
C2250 addersubtractor_0/XOR_1/NAND_3/a_6_n14# Gnd 0.14fF
C2251 addersubtractor_0/XOR_1/NAND_3/in2 Gnd 0.76fF
C2252 addersubtractor_0/XOR_1/NAND_3/w_32_0# Gnd 0.40fF
C2253 addersubtractor_0/XOR_1/NAND_3/w_0_0# Gnd 0.40fF
C2254 addersubtractor_0/XOR_1/NAND_2/a_6_n14# Gnd 0.14fF
C2255 addersubtractor_0/XOR_1/NAND_2/w_32_0# Gnd 0.40fF
C2256 addersubtractor_0/XOR_1/NAND_2/w_0_0# Gnd 0.40fF
C2257 addersubtractor_0/XOR_1/NAND_1/a_6_n14# Gnd 0.14fF
C2258 addersubtractor_0/XOR_1/NAND_3/in1 Gnd 0.78fF
C2259 addersubtractor_0/XOR_1/NAND_1/w_32_0# Gnd 0.40fF
C2260 addersubtractor_0/XOR_1/NAND_1/w_0_0# Gnd 0.40fF
C2261 addersubtractor_0/XOR_1/NAND_0/a_6_n14# Gnd 0.14fF
C2262 addersubtractor_0/XOR_1/NAND_2/in1 Gnd 0.97fF
C2263 addersubtractor_0/XOR_1/NAND_0/w_32_0# Gnd 0.40fF
C2264 addersubtractor_0/XOR_1/NAND_0/w_0_0# Gnd 0.40fF
C2265 addersubtractor_0/fulladder_3/XOR_1/NAND_3/a_6_n14# Gnd 0.14fF
C2266 adder3 Gnd 0.51fF
C2267 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 Gnd 0.76fF
C2268 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_32_0# Gnd 0.40fF
C2269 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_0_0# Gnd 0.40fF
C2270 addersubtractor_0/fulladder_3/XOR_1/NAND_2/a_6_n14# Gnd 0.14fF
C2271 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_32_0# Gnd 0.40fF
C2272 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_0_0# Gnd 0.40fF
C2273 addersubtractor_0/fulladder_3/XOR_1/NAND_1/a_6_n14# Gnd 0.14fF
C2274 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 Gnd 0.78fF
C2275 addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_32_0# Gnd 0.40fF
C2276 addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_0_0# Gnd 0.40fF
C2277 addersubtractor_0/fulladder_3/XOR_1/NAND_0/a_6_n14# Gnd 0.14fF
C2278 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 Gnd 0.97fF
C2279 addersubtractor_0/fulladder_2/C Gnd 1.24fF
C2280 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_32_0# Gnd 0.40fF
C2281 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_0_0# Gnd 0.40fF
C2282 addersubtractor_0/fulladder_3/OR_0/NOT_0/in Gnd 0.77fF
C2283 addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# Gnd 0.02fF
C2284 addersubtractor_0/fulladder_3/OR_0/in1 Gnd 0.40fF
C2285 addersubtractor_0/fulladder_3/OR_0/NOR_0/w_32_0# Gnd 0.40fF
C2286 addersubtractor_0/fulladder_3/OR_0/NOR_0/w_0_0# Gnd 0.40fF
C2287 AND_0/in1 Gnd 0.43fF
C2288 addersubtractor_0/fulladder_3/OR_0/NOT_0/w_0_0# Gnd 0.40fF
C2289 addersubtractor_0/fulladder_3/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C2290 addersubtractor_0/fulladder_3/XOR_1/in2 Gnd 2.44fF
C2291 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 Gnd 0.76fF
C2292 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C2293 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C2294 addersubtractor_0/fulladder_3/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C2295 addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C2296 addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C2297 addersubtractor_0/fulladder_3/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C2298 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 Gnd 0.78fF
C2299 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C2300 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C2301 addersubtractor_0/fulladder_3/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C2302 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 Gnd 0.97fF
C2303 addersubtractor_0/XOR_3/out Gnd 1.88fF
C2304 enableblock_0/B_out1 Gnd 2.66fF
C2305 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C2306 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C2307 addersubtractor_0/fulladder_3/AND_1/not_0/in Gnd 0.76fF
C2308 addersubtractor_0/fulladder_3/AND_1/not_0/w_0_0# Gnd 0.40fF
C2309 addersubtractor_0/fulladder_3/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2310 addersubtractor_0/fulladder_3/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2311 addersubtractor_0/fulladder_3/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2312 addersubtractor_0/fulladder_3/AND_0/not_0/in Gnd 0.76fF
C2313 addersubtractor_0/fulladder_3/OR_0/in2 Gnd 0.47fF
C2314 addersubtractor_0/fulladder_3/AND_0/not_0/w_0_0# Gnd 0.40fF
C2315 addersubtractor_0/fulladder_3/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2316 addersubtractor_0/fulladder_3/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2317 addersubtractor_0/fulladder_3/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2318 addersubtractor_0/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C2319 addersubtractor_0/XOR_0/NAND_3/in2 Gnd 0.76fF
C2320 addersubtractor_0/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C2321 addersubtractor_0/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C2322 addersubtractor_0/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C2323 addersubtractor_0/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C2324 addersubtractor_0/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C2325 addersubtractor_0/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C2326 addersubtractor_0/XOR_0/NAND_3/in1 Gnd 0.78fF
C2327 addersubtractor_0/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C2328 addersubtractor_0/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C2329 addersubtractor_0/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C2330 addersubtractor_0/XOR_0/NAND_2/in1 Gnd 0.97fF
C2331 S0 Gnd 10.27fF
C2332 addersubtractor_0/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C2333 addersubtractor_0/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C2334 addersubtractor_0/fulladder_2/XOR_1/NAND_3/a_6_n14# Gnd 0.14fF
C2335 adder2 Gnd 0.57fF
C2336 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 Gnd 0.76fF
C2337 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_32_0# Gnd 0.40fF
C2338 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_0_0# Gnd 0.40fF
C2339 addersubtractor_0/fulladder_2/XOR_1/NAND_2/a_6_n14# Gnd 0.14fF
C2340 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_32_0# Gnd 0.40fF
C2341 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_0_0# Gnd 0.40fF
C2342 addersubtractor_0/fulladder_2/XOR_1/NAND_1/a_6_n14# Gnd 0.14fF
C2343 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 Gnd 0.78fF
C2344 addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_32_0# Gnd 0.40fF
C2345 addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_0_0# Gnd 0.40fF
C2346 gnd Gnd 93.68fF
C2347 addersubtractor_0/fulladder_2/XOR_1/NAND_0/a_6_n14# Gnd 0.14fF
C2348 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 Gnd 0.97fF
C2349 addersubtractor_0/fulladder_1/C Gnd 1.25fF
C2350 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_32_0# Gnd 0.40fF
C2351 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_0_0# Gnd 0.40fF
C2352 addersubtractor_0/fulladder_2/OR_0/NOT_0/in Gnd 0.77fF
C2353 addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# Gnd 0.02fF
C2354 addersubtractor_0/fulladder_2/OR_0/in1 Gnd 0.40fF
C2355 addersubtractor_0/fulladder_2/OR_0/NOR_0/w_32_0# Gnd 0.40fF
C2356 addersubtractor_0/fulladder_2/OR_0/NOR_0/w_0_0# Gnd 0.40fF
C2357 addersubtractor_0/fulladder_2/OR_0/NOT_0/w_0_0# Gnd 0.40fF
C2358 addersubtractor_0/fulladder_2/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C2359 addersubtractor_0/fulladder_2/XOR_1/in2 Gnd 2.44fF
C2360 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 Gnd 0.76fF
C2361 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C2362 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C2363 addersubtractor_0/fulladder_2/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C2364 addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C2365 addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C2366 addersubtractor_0/fulladder_2/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C2367 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 Gnd 0.78fF
C2368 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C2369 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C2370 addersubtractor_0/fulladder_2/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C2371 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 Gnd 0.97fF
C2372 addersubtractor_0/XOR_2/out Gnd 1.88fF
C2373 enableblock_0/B_out3 Gnd 2.50fF
C2374 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C2375 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C2376 addersubtractor_0/fulladder_2/AND_1/not_0/in Gnd 0.76fF
C2377 addersubtractor_0/fulladder_2/AND_1/not_0/w_0_0# Gnd 0.40fF
C2378 addersubtractor_0/fulladder_2/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2379 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2380 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2381 addersubtractor_0/fulladder_2/AND_0/not_0/in Gnd 0.76fF
C2382 addersubtractor_0/fulladder_2/OR_0/in2 Gnd 0.47fF
C2383 addersubtractor_0/fulladder_2/AND_0/not_0/w_0_0# Gnd 0.40fF
C2384 addersubtractor_0/fulladder_2/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2385 addersubtractor_0/fulladder_2/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2386 addersubtractor_0/fulladder_2/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2387 addersubtractor_0/fulladder_1/XOR_1/NAND_3/a_6_n14# Gnd 0.14fF
C2388 adder1 Gnd 0.54fF
C2389 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 Gnd 0.76fF
C2390 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_32_0# Gnd 0.40fF
C2391 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_0_0# Gnd 0.40fF
C2392 addersubtractor_0/fulladder_1/XOR_1/NAND_2/a_6_n14# Gnd 0.14fF
C2393 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_32_0# Gnd 0.40fF
C2394 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_0_0# Gnd 0.40fF
C2395 addersubtractor_0/fulladder_1/XOR_1/NAND_1/a_6_n14# Gnd 0.14fF
C2396 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 Gnd 0.78fF
C2397 addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_32_0# Gnd 0.40fF
C2398 addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_0_0# Gnd 0.40fF
C2399 addersubtractor_0/fulladder_1/XOR_1/NAND_0/a_6_n14# Gnd 0.14fF
C2400 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 Gnd 0.97fF
C2401 addersubtractor_0/fulladder_0/C Gnd 1.23fF
C2402 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_32_0# Gnd 0.40fF
C2403 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_0_0# Gnd 0.40fF
C2404 addersubtractor_0/fulladder_1/OR_0/NOT_0/in Gnd 0.77fF
C2405 addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# Gnd 0.02fF
C2406 addersubtractor_0/fulladder_1/OR_0/in1 Gnd 0.40fF
C2407 addersubtractor_0/fulladder_1/OR_0/NOR_0/w_32_0# Gnd 0.40fF
C2408 addersubtractor_0/fulladder_1/OR_0/NOR_0/w_0_0# Gnd 0.40fF
C2409 addersubtractor_0/fulladder_1/OR_0/NOT_0/w_0_0# Gnd 0.40fF
C2410 addersubtractor_0/fulladder_1/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C2411 addersubtractor_0/fulladder_1/XOR_1/in2 Gnd 2.44fF
C2412 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 Gnd 0.76fF
C2413 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C2414 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C2415 addersubtractor_0/fulladder_1/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C2416 addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C2417 addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C2418 addersubtractor_0/fulladder_1/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C2419 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 Gnd 0.78fF
C2420 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C2421 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C2422 addersubtractor_0/fulladder_1/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C2423 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 Gnd 0.97fF
C2424 addersubtractor_0/XOR_1/out Gnd 1.88fF
C2425 enableblock_0/A_out1 Gnd 2.48fF
C2426 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C2427 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C2428 addersubtractor_0/fulladder_1/AND_1/not_0/in Gnd 0.76fF
C2429 addersubtractor_0/fulladder_1/AND_1/not_0/w_0_0# Gnd 0.40fF
C2430 addersubtractor_0/fulladder_1/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2431 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2432 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2433 addersubtractor_0/fulladder_1/AND_0/not_0/in Gnd 0.76fF
C2434 addersubtractor_0/fulladder_1/OR_0/in2 Gnd 0.47fF
C2435 addersubtractor_0/fulladder_1/AND_0/not_0/w_0_0# Gnd 0.40fF
C2436 addersubtractor_0/fulladder_1/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2437 addersubtractor_0/fulladder_1/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2438 addersubtractor_0/fulladder_1/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2439 addersubtractor_0/fulladder_0/XOR_1/NAND_3/a_6_n14# Gnd 0.14fF
C2440 adder0 Gnd 0.57fF
C2441 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 Gnd 0.76fF
C2442 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_32_0# Gnd 0.40fF
C2443 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_0_0# Gnd 0.40fF
C2444 addersubtractor_0/fulladder_0/XOR_1/NAND_2/a_6_n14# Gnd 0.14fF
C2445 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_32_0# Gnd 0.40fF
C2446 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_0_0# Gnd 0.40fF
C2447 addersubtractor_0/fulladder_0/XOR_1/NAND_1/a_6_n14# Gnd 0.14fF
C2448 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 Gnd 0.78fF
C2449 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_32_0# Gnd 0.40fF
C2450 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_0_0# Gnd 0.40fF
C2451 addersubtractor_0/fulladder_0/XOR_1/NAND_0/a_6_n14# Gnd 0.14fF
C2452 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 Gnd 0.97fF
C2453 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_32_0# Gnd 0.40fF
C2454 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_0_0# Gnd 0.40fF
C2455 addersubtractor_0/fulladder_0/OR_0/NOT_0/in Gnd 0.77fF
C2456 addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# Gnd 0.02fF
C2457 addersubtractor_0/fulladder_0/OR_0/in1 Gnd 0.40fF
C2458 addersubtractor_0/fulladder_0/OR_0/NOR_0/w_32_0# Gnd 0.40fF
C2459 addersubtractor_0/fulladder_0/OR_0/NOR_0/w_0_0# Gnd 0.40fF
C2460 addersubtractor_0/fulladder_0/OR_0/NOT_0/w_0_0# Gnd 0.40fF
C2461 vdd Gnd 29.45fF
C2462 addersubtractor_0/fulladder_0/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C2463 addersubtractor_0/fulladder_0/XOR_1/in2 Gnd 2.44fF
C2464 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 Gnd 0.76fF
C2465 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C2466 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C2467 addersubtractor_0/fulladder_0/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C2468 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C2469 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C2470 addersubtractor_0/fulladder_0/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C2471 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 Gnd 0.78fF
C2472 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C2473 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C2474 addersubtractor_0/fulladder_0/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C2475 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 Gnd 0.97fF
C2476 addersubtractor_0/XOR_0/out Gnd 1.87fF
C2477 enableblock_0/A_out3 Gnd 3.35fF
C2478 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C2479 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C2480 addersubtractor_0/fulladder_0/AND_1/not_0/in Gnd 0.76fF
C2481 addersubtractor_0/fulladder_0/AND_1/not_0/w_0_0# Gnd 0.40fF
C2482 addersubtractor_0/fulladder_0/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2483 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2484 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2485 addersubtractor_0/fulladder_0/AND_0/not_0/in Gnd 0.76fF
C2486 addersubtractor_0/fulladder_0/OR_0/in2 Gnd 0.47fF
C2487 addersubtractor_0/fulladder_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C2488 addersubtractor_0/fulladder_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2489 addersubtractor_0/fulladder_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2490 vdd Gnd 0.40fF


.tran 1n 400n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(node_A0) v(node_A1)+2 v(node_A2)+4 v(node_A3)+6 v(node_B0)+8 v(node_B1)+10 v(node_B2)+12 v(node_B3)+14
plot v(S0) v(S1)+2 v(adder0)+4 v(adder1)+6 v(adder2)+8 v(adder3)+10 v(carry)+12
plot v(S0) v(S1)+2 v(lesser)+4 v(equal)+6 v(greater)+8 
plot v(S0) v(S1)+2 v(and0)+4 v(and1)+6 v(and2)+8 v(and3)+10 
.end
.endc